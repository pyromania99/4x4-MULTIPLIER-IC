magic
tech scmos
timestamp 1668811232
<< nwell >>
rect -4671 1577 -4603 1597
rect -4586 1577 -4541 1597
rect -4671 1477 -4603 1497
rect -4586 1477 -4541 1497
rect -4290 1428 -4222 1448
rect -4003 1428 -3935 1448
rect -3658 1429 -3590 1449
rect -3343 1429 -3275 1449
rect -4671 1370 -4603 1390
rect -4586 1370 -4541 1390
rect -4371 1353 -4303 1373
rect -4204 1350 -4136 1370
rect -4084 1353 -4016 1373
rect -3917 1350 -3849 1370
rect -3739 1354 -3671 1374
rect -3572 1351 -3504 1371
rect -3424 1354 -3356 1374
rect -3257 1351 -3189 1371
rect -4671 1270 -4603 1290
rect -4586 1270 -4541 1290
rect -4290 1268 -4222 1288
rect -4003 1268 -3935 1288
rect -3658 1269 -3590 1289
rect -3343 1269 -3275 1289
rect -4671 1167 -4603 1187
rect -4586 1167 -4541 1187
rect -4367 1162 -4299 1182
rect -4282 1162 -4237 1182
rect -4080 1162 -4012 1182
rect -3995 1162 -3950 1182
rect -3933 1156 -3869 1177
rect -3860 1156 -3821 1177
rect -3735 1163 -3667 1183
rect -3650 1163 -3605 1183
rect -3420 1163 -3352 1183
rect -3335 1163 -3290 1183
rect -3273 1157 -3209 1178
rect -3200 1157 -3161 1178
rect -4671 1067 -4603 1087
rect -4586 1067 -4541 1087
rect -4290 1012 -4222 1032
rect -4003 1012 -3935 1032
rect -3657 1012 -3589 1032
rect -3375 1012 -3307 1032
rect -3048 1017 -2980 1037
rect -4671 960 -4603 980
rect -4586 960 -4541 980
rect -4371 937 -4303 957
rect -4204 934 -4136 954
rect -4084 937 -4016 957
rect -3917 934 -3849 954
rect -3738 937 -3670 957
rect -3571 934 -3503 954
rect -3456 937 -3388 957
rect -3289 934 -3221 954
rect -3129 942 -3061 962
rect -2962 939 -2894 959
rect -4671 860 -4603 880
rect -4586 860 -4541 880
rect -4290 852 -4222 872
rect -4003 852 -3935 872
rect -3657 852 -3589 872
rect -3375 852 -3307 872
rect -3048 857 -2980 877
rect -4672 745 -4604 765
rect -4587 745 -4542 765
rect -4367 746 -4299 766
rect -4282 746 -4237 766
rect -4080 746 -4012 766
rect -3995 746 -3950 766
rect -3933 740 -3869 761
rect -3860 740 -3821 761
rect -3734 746 -3666 766
rect -3649 746 -3604 766
rect -3452 746 -3384 766
rect -3367 746 -3322 766
rect -3305 740 -3241 761
rect -3232 740 -3193 761
rect -3125 751 -3057 771
rect -3040 751 -2995 771
rect -4672 645 -4604 665
rect -4587 645 -4542 665
rect -4672 538 -4604 558
rect -4587 538 -4542 558
rect -4290 554 -4222 574
rect -3991 554 -3923 574
rect -3676 554 -3608 574
rect -3347 560 -3279 580
rect -3032 560 -2964 580
rect -4371 479 -4303 499
rect -4204 476 -4136 496
rect -4072 479 -4004 499
rect -3905 476 -3837 496
rect -3757 479 -3689 499
rect -3590 476 -3522 496
rect -3428 485 -3360 505
rect -3261 482 -3193 502
rect -3113 485 -3045 505
rect -2946 482 -2878 502
rect -4672 438 -4604 458
rect -4587 438 -4542 458
rect -4290 394 -4222 414
rect -3991 394 -3923 414
rect -3676 394 -3608 414
rect -3347 400 -3279 420
rect -3032 400 -2964 420
rect -4672 335 -4604 355
rect -4587 335 -4542 355
rect -4367 288 -4299 308
rect -4282 288 -4237 308
rect -4068 288 -4000 308
rect -3983 288 -3938 308
rect -3753 288 -3685 308
rect -3668 288 -3623 308
rect -3424 294 -3356 314
rect -3339 294 -3294 314
rect -3109 294 -3041 314
rect -3024 294 -2979 314
rect -3606 262 -3542 283
rect -3533 262 -3494 283
rect -2962 268 -2898 289
rect -2889 268 -2850 289
rect -4672 235 -4604 255
rect -4587 235 -4542 255
rect -4290 180 -4222 200
rect -4672 128 -4604 148
rect -4587 128 -4542 148
rect -3959 147 -3891 167
rect -3644 147 -3576 167
rect -4371 105 -4303 125
rect -4204 102 -4136 122
rect -4040 72 -3972 92
rect -3873 69 -3805 89
rect -3725 72 -3657 92
rect -3558 69 -3490 89
rect -4672 28 -4604 48
rect -4587 28 -4542 48
rect -4290 20 -4222 40
rect -3959 -13 -3891 7
rect -3644 -13 -3576 7
rect -4367 -86 -4299 -66
rect -4282 -86 -4237 -66
rect -4036 -119 -3968 -99
rect -3951 -119 -3906 -99
rect -3721 -119 -3653 -99
rect -3636 -119 -3591 -99
rect -3574 -145 -3510 -124
rect -3501 -145 -3462 -124
rect -4290 -196 -4222 -176
rect -4371 -271 -4303 -251
rect -4204 -274 -4136 -254
rect -4290 -356 -4222 -336
rect -4367 -462 -4299 -442
rect -4282 -462 -4237 -442
<< ntransistor >>
rect -4656 1534 -4651 1543
rect -4628 1534 -4623 1543
rect -4571 1534 -4566 1543
rect -4656 1434 -4651 1443
rect -4628 1434 -4623 1443
rect -4571 1434 -4566 1443
rect -4275 1385 -4270 1394
rect -4247 1385 -4242 1394
rect -4656 1327 -4651 1336
rect -4628 1327 -4623 1336
rect -4571 1327 -4566 1336
rect -3988 1385 -3983 1394
rect -3960 1385 -3955 1394
rect -4356 1310 -4351 1319
rect -4328 1310 -4323 1319
rect -3643 1386 -3638 1395
rect -3615 1386 -3610 1395
rect -4189 1307 -4184 1316
rect -4161 1307 -4156 1316
rect -4069 1310 -4064 1319
rect -4041 1310 -4036 1319
rect -4656 1227 -4651 1236
rect -4628 1227 -4623 1236
rect -4571 1227 -4566 1236
rect -3328 1386 -3323 1395
rect -3300 1386 -3295 1395
rect -3902 1307 -3897 1316
rect -3874 1307 -3869 1316
rect -3724 1311 -3719 1320
rect -3696 1311 -3691 1320
rect -4275 1225 -4270 1234
rect -4247 1225 -4242 1234
rect -3557 1308 -3552 1317
rect -3529 1308 -3524 1317
rect -3409 1311 -3404 1320
rect -3381 1311 -3376 1320
rect -3988 1225 -3983 1234
rect -3960 1225 -3955 1234
rect -4656 1124 -4651 1133
rect -4628 1124 -4623 1133
rect -4571 1124 -4566 1133
rect -3242 1308 -3237 1317
rect -3214 1308 -3209 1317
rect -3643 1226 -3638 1235
rect -3615 1226 -3610 1235
rect -3328 1226 -3323 1235
rect -3300 1226 -3295 1235
rect -4352 1119 -4347 1128
rect -4324 1119 -4319 1128
rect -4267 1119 -4262 1128
rect -4065 1119 -4060 1128
rect -4037 1119 -4032 1128
rect -3980 1119 -3975 1128
rect -3919 1120 -3915 1125
rect -3892 1120 -3888 1125
rect -3844 1120 -3839 1125
rect -3720 1120 -3715 1129
rect -3692 1120 -3687 1129
rect -3635 1120 -3630 1129
rect -3405 1120 -3400 1129
rect -3377 1120 -3372 1129
rect -3320 1120 -3315 1129
rect -3259 1121 -3255 1126
rect -3232 1121 -3228 1126
rect -3184 1121 -3179 1126
rect -4656 1024 -4651 1033
rect -4628 1024 -4623 1033
rect -4571 1024 -4566 1033
rect -4275 969 -4270 978
rect -4247 969 -4242 978
rect -4656 917 -4651 926
rect -4628 917 -4623 926
rect -4571 917 -4566 926
rect -3988 969 -3983 978
rect -3960 969 -3955 978
rect -4356 894 -4351 903
rect -4328 894 -4323 903
rect -3642 969 -3637 978
rect -3614 969 -3609 978
rect -4189 891 -4184 900
rect -4161 891 -4156 900
rect -4069 894 -4064 903
rect -4041 894 -4036 903
rect -4656 817 -4651 826
rect -4628 817 -4623 826
rect -4571 817 -4566 826
rect -3360 969 -3355 978
rect -3332 969 -3327 978
rect -3902 891 -3897 900
rect -3874 891 -3869 900
rect -3723 894 -3718 903
rect -3695 894 -3690 903
rect -4275 809 -4270 818
rect -4247 809 -4242 818
rect -3033 974 -3028 983
rect -3005 974 -3000 983
rect -3556 891 -3551 900
rect -3528 891 -3523 900
rect -3441 894 -3436 903
rect -3413 894 -3408 903
rect -3988 809 -3983 818
rect -3960 809 -3955 818
rect -3274 891 -3269 900
rect -3246 891 -3241 900
rect -3114 899 -3109 908
rect -3086 899 -3081 908
rect -3642 809 -3637 818
rect -3614 809 -3609 818
rect -2947 896 -2942 905
rect -2919 896 -2914 905
rect -3360 809 -3355 818
rect -3332 809 -3327 818
rect -3033 814 -3028 823
rect -3005 814 -3000 823
rect -4657 702 -4652 711
rect -4629 702 -4624 711
rect -4572 702 -4567 711
rect -4352 703 -4347 712
rect -4324 703 -4319 712
rect -4267 703 -4262 712
rect -4065 703 -4060 712
rect -4037 703 -4032 712
rect -3980 703 -3975 712
rect -3919 704 -3915 709
rect -3892 704 -3888 709
rect -3844 704 -3839 709
rect -3719 703 -3714 712
rect -3691 703 -3686 712
rect -3634 703 -3629 712
rect -3437 703 -3432 712
rect -3409 703 -3404 712
rect -3352 703 -3347 712
rect -3291 704 -3287 709
rect -3264 704 -3260 709
rect -3216 704 -3211 709
rect -3110 708 -3105 717
rect -3082 708 -3077 717
rect -3025 708 -3020 717
rect -4657 602 -4652 611
rect -4629 602 -4624 611
rect -4572 602 -4567 611
rect -4657 495 -4652 504
rect -4629 495 -4624 504
rect -4572 495 -4567 504
rect -4275 511 -4270 520
rect -4247 511 -4242 520
rect -3976 511 -3971 520
rect -3948 511 -3943 520
rect -4356 436 -4351 445
rect -4328 436 -4323 445
rect -4657 395 -4652 404
rect -4629 395 -4624 404
rect -4572 395 -4567 404
rect -3661 511 -3656 520
rect -3633 511 -3628 520
rect -4189 433 -4184 442
rect -4161 433 -4156 442
rect -4057 436 -4052 445
rect -4029 436 -4024 445
rect -3332 517 -3327 526
rect -3304 517 -3299 526
rect -3890 433 -3885 442
rect -3862 433 -3857 442
rect -3742 436 -3737 445
rect -3714 436 -3709 445
rect -4275 351 -4270 360
rect -4247 351 -4242 360
rect -3017 517 -3012 526
rect -2989 517 -2984 526
rect -3413 442 -3408 451
rect -3385 442 -3380 451
rect -3575 433 -3570 442
rect -3547 433 -3542 442
rect -3976 351 -3971 360
rect -3948 351 -3943 360
rect -3246 439 -3241 448
rect -3218 439 -3213 448
rect -3098 442 -3093 451
rect -3070 442 -3065 451
rect -3661 351 -3656 360
rect -3633 351 -3628 360
rect -2931 439 -2926 448
rect -2903 439 -2898 448
rect -3332 357 -3327 366
rect -3304 357 -3299 366
rect -3017 357 -3012 366
rect -2989 357 -2984 366
rect -4657 292 -4652 301
rect -4629 292 -4624 301
rect -4572 292 -4567 301
rect -4352 245 -4347 254
rect -4324 245 -4319 254
rect -4267 245 -4262 254
rect -4053 245 -4048 254
rect -4025 245 -4020 254
rect -3968 245 -3963 254
rect -3738 245 -3733 254
rect -3710 245 -3705 254
rect -3653 245 -3648 254
rect -3409 251 -3404 260
rect -3381 251 -3376 260
rect -3324 251 -3319 260
rect -3094 251 -3089 260
rect -3066 251 -3061 260
rect -3009 251 -3004 260
rect -3592 226 -3588 231
rect -3565 226 -3561 231
rect -3517 226 -3512 231
rect -2948 232 -2944 237
rect -2921 232 -2917 237
rect -2873 232 -2868 237
rect -4657 192 -4652 201
rect -4629 192 -4624 201
rect -4572 192 -4567 201
rect -4275 137 -4270 146
rect -4247 137 -4242 146
rect -4657 85 -4652 94
rect -4629 85 -4624 94
rect -4572 85 -4567 94
rect -4356 62 -4351 71
rect -4328 62 -4323 71
rect -3944 104 -3939 113
rect -3916 104 -3911 113
rect -4189 59 -4184 68
rect -4161 59 -4156 68
rect -4657 -15 -4652 -6
rect -4629 -15 -4624 -6
rect -4572 -15 -4567 -6
rect -3629 104 -3624 113
rect -3601 104 -3596 113
rect -4025 29 -4020 38
rect -3997 29 -3992 38
rect -4275 -23 -4270 -14
rect -4247 -23 -4242 -14
rect -3858 26 -3853 35
rect -3830 26 -3825 35
rect -3710 29 -3705 38
rect -3682 29 -3677 38
rect -3543 26 -3538 35
rect -3515 26 -3510 35
rect -3944 -56 -3939 -47
rect -3916 -56 -3911 -47
rect -3629 -56 -3624 -47
rect -3601 -56 -3596 -47
rect -4352 -129 -4347 -120
rect -4324 -129 -4319 -120
rect -4267 -129 -4262 -120
rect -4021 -162 -4016 -153
rect -3993 -162 -3988 -153
rect -3936 -162 -3931 -153
rect -3706 -162 -3701 -153
rect -3678 -162 -3673 -153
rect -3621 -162 -3616 -153
rect -3560 -181 -3556 -176
rect -3533 -181 -3529 -176
rect -3485 -181 -3480 -176
rect -4275 -239 -4270 -230
rect -4247 -239 -4242 -230
rect -4356 -314 -4351 -305
rect -4328 -314 -4323 -305
rect -4189 -317 -4184 -308
rect -4161 -317 -4156 -308
rect -4275 -399 -4270 -390
rect -4247 -399 -4242 -390
rect -4352 -505 -4347 -496
rect -4324 -505 -4319 -496
rect -4267 -505 -4262 -496
<< ptransistor >>
rect -4656 1583 -4651 1591
rect -4628 1583 -4623 1591
rect -4571 1583 -4566 1591
rect -4656 1483 -4651 1491
rect -4628 1483 -4623 1491
rect -4571 1483 -4566 1491
rect -4275 1434 -4270 1442
rect -4247 1434 -4242 1442
rect -3988 1434 -3983 1442
rect -3960 1434 -3955 1442
rect -3643 1435 -3638 1443
rect -3615 1435 -3610 1443
rect -3328 1435 -3323 1443
rect -3300 1435 -3295 1443
rect -4656 1376 -4651 1384
rect -4628 1376 -4623 1384
rect -4571 1376 -4566 1384
rect -4356 1359 -4351 1367
rect -4328 1359 -4323 1367
rect -4189 1356 -4184 1364
rect -4161 1356 -4156 1364
rect -4069 1359 -4064 1367
rect -4041 1359 -4036 1367
rect -4656 1276 -4651 1284
rect -4628 1276 -4623 1284
rect -4571 1276 -4566 1284
rect -3902 1356 -3897 1364
rect -3874 1356 -3869 1364
rect -3724 1360 -3719 1368
rect -3696 1360 -3691 1368
rect -4275 1274 -4270 1282
rect -4247 1274 -4242 1282
rect -3557 1357 -3552 1365
rect -3529 1357 -3524 1365
rect -3409 1360 -3404 1368
rect -3381 1360 -3376 1368
rect -3988 1274 -3983 1282
rect -3960 1274 -3955 1282
rect -3242 1357 -3237 1365
rect -3214 1357 -3209 1365
rect -3643 1275 -3638 1283
rect -3615 1275 -3610 1283
rect -4656 1173 -4651 1181
rect -4628 1173 -4623 1181
rect -4571 1173 -4566 1181
rect -4352 1168 -4347 1176
rect -4324 1168 -4319 1176
rect -4267 1168 -4262 1176
rect -4065 1168 -4060 1176
rect -4037 1168 -4032 1176
rect -3980 1168 -3975 1176
rect -3328 1275 -3323 1283
rect -3300 1275 -3295 1283
rect -3919 1162 -3915 1171
rect -3892 1162 -3888 1171
rect -3844 1162 -3839 1171
rect -3720 1169 -3715 1177
rect -3692 1169 -3687 1177
rect -3635 1169 -3630 1177
rect -3405 1169 -3400 1177
rect -3377 1169 -3372 1177
rect -3320 1169 -3315 1177
rect -3259 1163 -3255 1172
rect -3232 1163 -3228 1172
rect -3184 1163 -3179 1172
rect -4656 1073 -4651 1081
rect -4628 1073 -4623 1081
rect -4571 1073 -4566 1081
rect -4275 1018 -4270 1026
rect -4247 1018 -4242 1026
rect -3988 1018 -3983 1026
rect -3960 1018 -3955 1026
rect -3642 1018 -3637 1026
rect -3614 1018 -3609 1026
rect -3360 1018 -3355 1026
rect -3332 1018 -3327 1026
rect -3033 1023 -3028 1031
rect -3005 1023 -3000 1031
rect -4656 966 -4651 974
rect -4628 966 -4623 974
rect -4571 966 -4566 974
rect -4356 943 -4351 951
rect -4328 943 -4323 951
rect -4189 940 -4184 948
rect -4161 940 -4156 948
rect -4069 943 -4064 951
rect -4041 943 -4036 951
rect -4656 866 -4651 874
rect -4628 866 -4623 874
rect -4571 866 -4566 874
rect -3902 940 -3897 948
rect -3874 940 -3869 948
rect -3723 943 -3718 951
rect -3695 943 -3690 951
rect -4275 858 -4270 866
rect -4247 858 -4242 866
rect -3556 940 -3551 948
rect -3528 940 -3523 948
rect -3441 943 -3436 951
rect -3413 943 -3408 951
rect -3988 858 -3983 866
rect -3960 858 -3955 866
rect -3114 948 -3109 956
rect -3086 948 -3081 956
rect -3274 940 -3269 948
rect -3246 940 -3241 948
rect -3642 858 -3637 866
rect -3614 858 -3609 866
rect -4657 751 -4652 759
rect -4629 751 -4624 759
rect -4572 751 -4567 759
rect -4352 752 -4347 760
rect -4324 752 -4319 760
rect -4267 752 -4262 760
rect -4065 752 -4060 760
rect -4037 752 -4032 760
rect -3980 752 -3975 760
rect -2947 945 -2942 953
rect -2919 945 -2914 953
rect -3360 858 -3355 866
rect -3332 858 -3327 866
rect -3033 863 -3028 871
rect -3005 863 -3000 871
rect -3919 746 -3915 755
rect -3892 746 -3888 755
rect -3844 746 -3839 755
rect -3719 752 -3714 760
rect -3691 752 -3686 760
rect -3634 752 -3629 760
rect -3437 752 -3432 760
rect -3409 752 -3404 760
rect -3352 752 -3347 760
rect -3110 757 -3105 765
rect -3082 757 -3077 765
rect -3025 757 -3020 765
rect -3291 746 -3287 755
rect -3264 746 -3260 755
rect -3216 746 -3211 755
rect -4657 651 -4652 659
rect -4629 651 -4624 659
rect -4572 651 -4567 659
rect -4275 560 -4270 568
rect -4247 560 -4242 568
rect -3976 560 -3971 568
rect -3948 560 -3943 568
rect -3661 560 -3656 568
rect -3633 560 -3628 568
rect -3332 566 -3327 574
rect -3304 566 -3299 574
rect -3017 566 -3012 574
rect -2989 566 -2984 574
rect -4657 544 -4652 552
rect -4629 544 -4624 552
rect -4572 544 -4567 552
rect -4356 485 -4351 493
rect -4328 485 -4323 493
rect -4657 444 -4652 452
rect -4629 444 -4624 452
rect -4572 444 -4567 452
rect -4189 482 -4184 490
rect -4161 482 -4156 490
rect -4057 485 -4052 493
rect -4029 485 -4024 493
rect -3890 482 -3885 490
rect -3862 482 -3857 490
rect -3742 485 -3737 493
rect -3714 485 -3709 493
rect -4275 400 -4270 408
rect -4247 400 -4242 408
rect -4657 341 -4652 349
rect -4629 341 -4624 349
rect -4572 341 -4567 349
rect -3413 491 -3408 499
rect -3385 491 -3380 499
rect -3575 482 -3570 490
rect -3547 482 -3542 490
rect -3976 400 -3971 408
rect -3948 400 -3943 408
rect -3246 488 -3241 496
rect -3218 488 -3213 496
rect -3098 491 -3093 499
rect -3070 491 -3065 499
rect -3661 400 -3656 408
rect -3633 400 -3628 408
rect -2931 488 -2926 496
rect -2903 488 -2898 496
rect -3332 406 -3327 414
rect -3304 406 -3299 414
rect -3017 406 -3012 414
rect -2989 406 -2984 414
rect -4352 294 -4347 302
rect -4324 294 -4319 302
rect -4267 294 -4262 302
rect -4053 294 -4048 302
rect -4025 294 -4020 302
rect -3968 294 -3963 302
rect -3738 294 -3733 302
rect -3710 294 -3705 302
rect -3653 294 -3648 302
rect -3409 300 -3404 308
rect -3381 300 -3376 308
rect -3324 300 -3319 308
rect -3094 300 -3089 308
rect -3066 300 -3061 308
rect -3009 300 -3004 308
rect -3592 268 -3588 277
rect -3565 268 -3561 277
rect -3517 268 -3512 277
rect -4657 241 -4652 249
rect -4629 241 -4624 249
rect -4572 241 -4567 249
rect -2948 274 -2944 283
rect -2921 274 -2917 283
rect -2873 274 -2868 283
rect -4275 186 -4270 194
rect -4247 186 -4242 194
rect -4657 134 -4652 142
rect -4629 134 -4624 142
rect -4572 134 -4567 142
rect -4356 111 -4351 119
rect -4328 111 -4323 119
rect -3944 153 -3939 161
rect -3916 153 -3911 161
rect -3629 153 -3624 161
rect -3601 153 -3596 161
rect -4189 108 -4184 116
rect -4161 108 -4156 116
rect -4657 34 -4652 42
rect -4629 34 -4624 42
rect -4572 34 -4567 42
rect -4025 78 -4020 86
rect -3997 78 -3992 86
rect -4275 26 -4270 34
rect -4247 26 -4242 34
rect -3858 75 -3853 83
rect -3830 75 -3825 83
rect -3710 78 -3705 86
rect -3682 78 -3677 86
rect -3543 75 -3538 83
rect -3515 75 -3510 83
rect -3944 -7 -3939 1
rect -3916 -7 -3911 1
rect -4352 -80 -4347 -72
rect -4324 -80 -4319 -72
rect -4267 -80 -4262 -72
rect -3629 -7 -3624 1
rect -3601 -7 -3596 1
rect -4021 -113 -4016 -105
rect -3993 -113 -3988 -105
rect -3936 -113 -3931 -105
rect -3706 -113 -3701 -105
rect -3678 -113 -3673 -105
rect -3621 -113 -3616 -105
rect -3560 -139 -3556 -130
rect -3533 -139 -3529 -130
rect -3485 -139 -3480 -130
rect -4275 -190 -4270 -182
rect -4247 -190 -4242 -182
rect -4356 -265 -4351 -257
rect -4328 -265 -4323 -257
rect -4189 -268 -4184 -260
rect -4161 -268 -4156 -260
rect -4275 -350 -4270 -342
rect -4247 -350 -4242 -342
rect -4352 -456 -4347 -448
rect -4324 -456 -4319 -448
rect -4267 -456 -4262 -448
<< ndiffusion >>
rect -4662 1534 -4656 1543
rect -4651 1534 -4628 1543
rect -4623 1534 -4616 1543
rect -4579 1534 -4571 1543
rect -4566 1534 -4558 1543
rect -4662 1434 -4656 1443
rect -4651 1434 -4628 1443
rect -4623 1434 -4616 1443
rect -4579 1434 -4571 1443
rect -4566 1434 -4558 1443
rect -4281 1385 -4275 1394
rect -4270 1385 -4247 1394
rect -4242 1385 -4235 1394
rect -4662 1327 -4656 1336
rect -4651 1327 -4628 1336
rect -4623 1327 -4616 1336
rect -4579 1327 -4571 1336
rect -4566 1327 -4558 1336
rect -3994 1385 -3988 1394
rect -3983 1385 -3960 1394
rect -3955 1385 -3948 1394
rect -4362 1310 -4356 1319
rect -4351 1310 -4328 1319
rect -4323 1310 -4316 1319
rect -3649 1386 -3643 1395
rect -3638 1386 -3615 1395
rect -3610 1386 -3603 1395
rect -4195 1307 -4189 1316
rect -4184 1307 -4161 1316
rect -4156 1307 -4149 1316
rect -4075 1310 -4069 1319
rect -4064 1310 -4041 1319
rect -4036 1310 -4029 1319
rect -4662 1227 -4656 1236
rect -4651 1227 -4628 1236
rect -4623 1227 -4616 1236
rect -4579 1227 -4571 1236
rect -4566 1227 -4558 1236
rect -3334 1386 -3328 1395
rect -3323 1386 -3300 1395
rect -3295 1386 -3288 1395
rect -3908 1307 -3902 1316
rect -3897 1307 -3874 1316
rect -3869 1307 -3862 1316
rect -3730 1311 -3724 1320
rect -3719 1311 -3696 1320
rect -3691 1311 -3684 1320
rect -4281 1225 -4275 1234
rect -4270 1225 -4247 1234
rect -4242 1225 -4235 1234
rect -3563 1308 -3557 1317
rect -3552 1308 -3529 1317
rect -3524 1308 -3517 1317
rect -3415 1311 -3409 1320
rect -3404 1311 -3381 1320
rect -3376 1311 -3369 1320
rect -3994 1225 -3988 1234
rect -3983 1225 -3960 1234
rect -3955 1225 -3948 1234
rect -4662 1124 -4656 1133
rect -4651 1124 -4628 1133
rect -4623 1124 -4616 1133
rect -4579 1124 -4571 1133
rect -4566 1124 -4558 1133
rect -3248 1308 -3242 1317
rect -3237 1308 -3214 1317
rect -3209 1308 -3202 1317
rect -3649 1226 -3643 1235
rect -3638 1226 -3615 1235
rect -3610 1226 -3603 1235
rect -3334 1226 -3328 1235
rect -3323 1226 -3300 1235
rect -3295 1226 -3288 1235
rect -4358 1119 -4352 1128
rect -4347 1119 -4324 1128
rect -4319 1119 -4312 1128
rect -4275 1119 -4267 1128
rect -4262 1119 -4254 1128
rect -4071 1119 -4065 1128
rect -4060 1119 -4037 1128
rect -4032 1119 -4025 1128
rect -3988 1119 -3980 1128
rect -3975 1119 -3967 1128
rect -3923 1120 -3919 1125
rect -3915 1120 -3908 1125
rect -3902 1120 -3892 1125
rect -3888 1120 -3882 1125
rect -3853 1120 -3844 1125
rect -3839 1120 -3833 1125
rect -3726 1120 -3720 1129
rect -3715 1120 -3692 1129
rect -3687 1120 -3680 1129
rect -3643 1120 -3635 1129
rect -3630 1120 -3622 1129
rect -3411 1120 -3405 1129
rect -3400 1120 -3377 1129
rect -3372 1120 -3365 1129
rect -3328 1120 -3320 1129
rect -3315 1120 -3307 1129
rect -3263 1121 -3259 1126
rect -3255 1121 -3248 1126
rect -3242 1121 -3232 1126
rect -3228 1121 -3222 1126
rect -3193 1121 -3184 1126
rect -3179 1121 -3173 1126
rect -4662 1024 -4656 1033
rect -4651 1024 -4628 1033
rect -4623 1024 -4616 1033
rect -4579 1024 -4571 1033
rect -4566 1024 -4558 1033
rect -4281 969 -4275 978
rect -4270 969 -4247 978
rect -4242 969 -4235 978
rect -4662 917 -4656 926
rect -4651 917 -4628 926
rect -4623 917 -4616 926
rect -4579 917 -4571 926
rect -4566 917 -4558 926
rect -3994 969 -3988 978
rect -3983 969 -3960 978
rect -3955 969 -3948 978
rect -4362 894 -4356 903
rect -4351 894 -4328 903
rect -4323 894 -4316 903
rect -3648 969 -3642 978
rect -3637 969 -3614 978
rect -3609 969 -3602 978
rect -4195 891 -4189 900
rect -4184 891 -4161 900
rect -4156 891 -4149 900
rect -4075 894 -4069 903
rect -4064 894 -4041 903
rect -4036 894 -4029 903
rect -4662 817 -4656 826
rect -4651 817 -4628 826
rect -4623 817 -4616 826
rect -4579 817 -4571 826
rect -4566 817 -4558 826
rect -3366 969 -3360 978
rect -3355 969 -3332 978
rect -3327 969 -3320 978
rect -3908 891 -3902 900
rect -3897 891 -3874 900
rect -3869 891 -3862 900
rect -3729 894 -3723 903
rect -3718 894 -3695 903
rect -3690 894 -3683 903
rect -4281 809 -4275 818
rect -4270 809 -4247 818
rect -4242 809 -4235 818
rect -3039 974 -3033 983
rect -3028 974 -3005 983
rect -3000 974 -2993 983
rect -3562 891 -3556 900
rect -3551 891 -3528 900
rect -3523 891 -3516 900
rect -3447 894 -3441 903
rect -3436 894 -3413 903
rect -3408 894 -3401 903
rect -3994 809 -3988 818
rect -3983 809 -3960 818
rect -3955 809 -3948 818
rect -3280 891 -3274 900
rect -3269 891 -3246 900
rect -3241 891 -3234 900
rect -3120 899 -3114 908
rect -3109 899 -3086 908
rect -3081 899 -3074 908
rect -3648 809 -3642 818
rect -3637 809 -3614 818
rect -3609 809 -3602 818
rect -2953 896 -2947 905
rect -2942 896 -2919 905
rect -2914 896 -2907 905
rect -3366 809 -3360 818
rect -3355 809 -3332 818
rect -3327 809 -3320 818
rect -3039 814 -3033 823
rect -3028 814 -3005 823
rect -3000 814 -2993 823
rect -4663 702 -4657 711
rect -4652 702 -4629 711
rect -4624 702 -4617 711
rect -4580 702 -4572 711
rect -4567 702 -4559 711
rect -4358 703 -4352 712
rect -4347 703 -4324 712
rect -4319 703 -4312 712
rect -4275 703 -4267 712
rect -4262 703 -4254 712
rect -4071 703 -4065 712
rect -4060 703 -4037 712
rect -4032 703 -4025 712
rect -3988 703 -3980 712
rect -3975 703 -3967 712
rect -3923 704 -3919 709
rect -3915 704 -3908 709
rect -3902 704 -3892 709
rect -3888 704 -3882 709
rect -3853 704 -3844 709
rect -3839 704 -3833 709
rect -3725 703 -3719 712
rect -3714 703 -3691 712
rect -3686 703 -3679 712
rect -3642 703 -3634 712
rect -3629 703 -3621 712
rect -3443 703 -3437 712
rect -3432 703 -3409 712
rect -3404 703 -3397 712
rect -3360 703 -3352 712
rect -3347 703 -3339 712
rect -3295 704 -3291 709
rect -3287 704 -3280 709
rect -3274 704 -3264 709
rect -3260 704 -3254 709
rect -3225 704 -3216 709
rect -3211 704 -3205 709
rect -3116 708 -3110 717
rect -3105 708 -3082 717
rect -3077 708 -3070 717
rect -3033 708 -3025 717
rect -3020 708 -3012 717
rect -4663 602 -4657 611
rect -4652 602 -4629 611
rect -4624 602 -4617 611
rect -4580 602 -4572 611
rect -4567 602 -4559 611
rect -4663 495 -4657 504
rect -4652 495 -4629 504
rect -4624 495 -4617 504
rect -4580 495 -4572 504
rect -4567 495 -4559 504
rect -4281 511 -4275 520
rect -4270 511 -4247 520
rect -4242 511 -4235 520
rect -3982 511 -3976 520
rect -3971 511 -3948 520
rect -3943 511 -3936 520
rect -4362 436 -4356 445
rect -4351 436 -4328 445
rect -4323 436 -4316 445
rect -4663 395 -4657 404
rect -4652 395 -4629 404
rect -4624 395 -4617 404
rect -4580 395 -4572 404
rect -4567 395 -4559 404
rect -3667 511 -3661 520
rect -3656 511 -3633 520
rect -3628 511 -3621 520
rect -4195 433 -4189 442
rect -4184 433 -4161 442
rect -4156 433 -4149 442
rect -4063 436 -4057 445
rect -4052 436 -4029 445
rect -4024 436 -4017 445
rect -3338 517 -3332 526
rect -3327 517 -3304 526
rect -3299 517 -3292 526
rect -3896 433 -3890 442
rect -3885 433 -3862 442
rect -3857 433 -3850 442
rect -3748 436 -3742 445
rect -3737 436 -3714 445
rect -3709 436 -3702 445
rect -4281 351 -4275 360
rect -4270 351 -4247 360
rect -4242 351 -4235 360
rect -3023 517 -3017 526
rect -3012 517 -2989 526
rect -2984 517 -2977 526
rect -3419 442 -3413 451
rect -3408 442 -3385 451
rect -3380 442 -3373 451
rect -3581 433 -3575 442
rect -3570 433 -3547 442
rect -3542 433 -3535 442
rect -3982 351 -3976 360
rect -3971 351 -3948 360
rect -3943 351 -3936 360
rect -3252 439 -3246 448
rect -3241 439 -3218 448
rect -3213 439 -3206 448
rect -3104 442 -3098 451
rect -3093 442 -3070 451
rect -3065 442 -3058 451
rect -3667 351 -3661 360
rect -3656 351 -3633 360
rect -3628 351 -3621 360
rect -2937 439 -2931 448
rect -2926 439 -2903 448
rect -2898 439 -2891 448
rect -3338 357 -3332 366
rect -3327 357 -3304 366
rect -3299 357 -3292 366
rect -3023 357 -3017 366
rect -3012 357 -2989 366
rect -2984 357 -2977 366
rect -4663 292 -4657 301
rect -4652 292 -4629 301
rect -4624 292 -4617 301
rect -4580 292 -4572 301
rect -4567 292 -4559 301
rect -4358 245 -4352 254
rect -4347 245 -4324 254
rect -4319 245 -4312 254
rect -4275 245 -4267 254
rect -4262 245 -4254 254
rect -4059 245 -4053 254
rect -4048 245 -4025 254
rect -4020 245 -4013 254
rect -3976 245 -3968 254
rect -3963 245 -3955 254
rect -3744 245 -3738 254
rect -3733 245 -3710 254
rect -3705 245 -3698 254
rect -3661 245 -3653 254
rect -3648 245 -3640 254
rect -3415 251 -3409 260
rect -3404 251 -3381 260
rect -3376 251 -3369 260
rect -3332 251 -3324 260
rect -3319 251 -3311 260
rect -3100 251 -3094 260
rect -3089 251 -3066 260
rect -3061 251 -3054 260
rect -3017 251 -3009 260
rect -3004 251 -2996 260
rect -3596 226 -3592 231
rect -3588 226 -3581 231
rect -3575 226 -3565 231
rect -3561 226 -3555 231
rect -3526 226 -3517 231
rect -3512 226 -3506 231
rect -2952 232 -2948 237
rect -2944 232 -2937 237
rect -2931 232 -2921 237
rect -2917 232 -2911 237
rect -2882 232 -2873 237
rect -2868 232 -2862 237
rect -4663 192 -4657 201
rect -4652 192 -4629 201
rect -4624 192 -4617 201
rect -4580 192 -4572 201
rect -4567 192 -4559 201
rect -4281 137 -4275 146
rect -4270 137 -4247 146
rect -4242 137 -4235 146
rect -4663 85 -4657 94
rect -4652 85 -4629 94
rect -4624 85 -4617 94
rect -4580 85 -4572 94
rect -4567 85 -4559 94
rect -4362 62 -4356 71
rect -4351 62 -4328 71
rect -4323 62 -4316 71
rect -3950 104 -3944 113
rect -3939 104 -3916 113
rect -3911 104 -3904 113
rect -4195 59 -4189 68
rect -4184 59 -4161 68
rect -4156 59 -4149 68
rect -4663 -15 -4657 -6
rect -4652 -15 -4629 -6
rect -4624 -15 -4617 -6
rect -4580 -15 -4572 -6
rect -4567 -15 -4559 -6
rect -3635 104 -3629 113
rect -3624 104 -3601 113
rect -3596 104 -3589 113
rect -4031 29 -4025 38
rect -4020 29 -3997 38
rect -3992 29 -3985 38
rect -4281 -23 -4275 -14
rect -4270 -23 -4247 -14
rect -4242 -23 -4235 -14
rect -3864 26 -3858 35
rect -3853 26 -3830 35
rect -3825 26 -3818 35
rect -3716 29 -3710 38
rect -3705 29 -3682 38
rect -3677 29 -3670 38
rect -3549 26 -3543 35
rect -3538 26 -3515 35
rect -3510 26 -3503 35
rect -3950 -56 -3944 -47
rect -3939 -56 -3916 -47
rect -3911 -56 -3904 -47
rect -3635 -56 -3629 -47
rect -3624 -56 -3601 -47
rect -3596 -56 -3589 -47
rect -4358 -129 -4352 -120
rect -4347 -129 -4324 -120
rect -4319 -129 -4312 -120
rect -4275 -129 -4267 -120
rect -4262 -129 -4254 -120
rect -4027 -162 -4021 -153
rect -4016 -162 -3993 -153
rect -3988 -162 -3981 -153
rect -3944 -162 -3936 -153
rect -3931 -162 -3923 -153
rect -3712 -162 -3706 -153
rect -3701 -162 -3678 -153
rect -3673 -162 -3666 -153
rect -3629 -162 -3621 -153
rect -3616 -162 -3608 -153
rect -3564 -181 -3560 -176
rect -3556 -181 -3549 -176
rect -3543 -181 -3533 -176
rect -3529 -181 -3523 -176
rect -3494 -181 -3485 -176
rect -3480 -181 -3474 -176
rect -4281 -239 -4275 -230
rect -4270 -239 -4247 -230
rect -4242 -239 -4235 -230
rect -4362 -314 -4356 -305
rect -4351 -314 -4328 -305
rect -4323 -314 -4316 -305
rect -4195 -317 -4189 -308
rect -4184 -317 -4161 -308
rect -4156 -317 -4149 -308
rect -4281 -399 -4275 -390
rect -4270 -399 -4247 -390
rect -4242 -399 -4235 -390
rect -4358 -505 -4352 -496
rect -4347 -505 -4324 -496
rect -4319 -505 -4312 -496
rect -4275 -505 -4267 -496
rect -4262 -505 -4254 -496
<< pdiffusion >>
rect -4658 1583 -4656 1591
rect -4651 1583 -4643 1591
rect -4636 1583 -4628 1591
rect -4623 1583 -4616 1591
rect -4573 1583 -4571 1591
rect -4566 1583 -4558 1591
rect -4551 1583 -4549 1591
rect -4658 1483 -4656 1491
rect -4651 1483 -4643 1491
rect -4636 1483 -4628 1491
rect -4623 1483 -4616 1491
rect -4573 1483 -4571 1491
rect -4566 1483 -4558 1491
rect -4551 1483 -4549 1491
rect -4277 1434 -4275 1442
rect -4270 1434 -4262 1442
rect -4255 1434 -4247 1442
rect -4242 1434 -4235 1442
rect -3990 1434 -3988 1442
rect -3983 1434 -3975 1442
rect -3968 1434 -3960 1442
rect -3955 1434 -3948 1442
rect -3645 1435 -3643 1443
rect -3638 1435 -3630 1443
rect -3623 1435 -3615 1443
rect -3610 1435 -3603 1443
rect -3330 1435 -3328 1443
rect -3323 1435 -3315 1443
rect -3308 1435 -3300 1443
rect -3295 1435 -3288 1443
rect -4658 1376 -4656 1384
rect -4651 1376 -4643 1384
rect -4636 1376 -4628 1384
rect -4623 1376 -4616 1384
rect -4573 1376 -4571 1384
rect -4566 1376 -4558 1384
rect -4551 1376 -4549 1384
rect -4358 1359 -4356 1367
rect -4351 1359 -4343 1367
rect -4336 1359 -4328 1367
rect -4323 1359 -4316 1367
rect -4191 1356 -4189 1364
rect -4184 1356 -4176 1364
rect -4169 1356 -4161 1364
rect -4156 1356 -4149 1364
rect -4071 1359 -4069 1367
rect -4064 1359 -4056 1367
rect -4049 1359 -4041 1367
rect -4036 1359 -4029 1367
rect -4658 1276 -4656 1284
rect -4651 1276 -4643 1284
rect -4636 1276 -4628 1284
rect -4623 1276 -4616 1284
rect -4573 1276 -4571 1284
rect -4566 1276 -4558 1284
rect -4551 1276 -4549 1284
rect -3904 1356 -3902 1364
rect -3897 1356 -3889 1364
rect -3882 1356 -3874 1364
rect -3869 1356 -3862 1364
rect -3726 1360 -3724 1368
rect -3719 1360 -3711 1368
rect -3704 1360 -3696 1368
rect -3691 1360 -3684 1368
rect -4277 1274 -4275 1282
rect -4270 1274 -4262 1282
rect -4255 1274 -4247 1282
rect -4242 1274 -4235 1282
rect -3559 1357 -3557 1365
rect -3552 1357 -3544 1365
rect -3537 1357 -3529 1365
rect -3524 1357 -3517 1365
rect -3411 1360 -3409 1368
rect -3404 1360 -3396 1368
rect -3389 1360 -3381 1368
rect -3376 1360 -3369 1368
rect -3990 1274 -3988 1282
rect -3983 1274 -3975 1282
rect -3968 1274 -3960 1282
rect -3955 1274 -3948 1282
rect -3244 1357 -3242 1365
rect -3237 1357 -3229 1365
rect -3222 1357 -3214 1365
rect -3209 1357 -3202 1365
rect -3645 1275 -3643 1283
rect -3638 1275 -3630 1283
rect -3623 1275 -3615 1283
rect -3610 1275 -3603 1283
rect -4658 1173 -4656 1181
rect -4651 1173 -4643 1181
rect -4636 1173 -4628 1181
rect -4623 1173 -4616 1181
rect -4573 1173 -4571 1181
rect -4566 1173 -4558 1181
rect -4551 1173 -4549 1181
rect -4354 1168 -4352 1176
rect -4347 1168 -4339 1176
rect -4332 1168 -4324 1176
rect -4319 1168 -4312 1176
rect -4269 1168 -4267 1176
rect -4262 1168 -4254 1176
rect -4247 1168 -4245 1176
rect -4067 1168 -4065 1176
rect -4060 1168 -4052 1176
rect -4045 1168 -4037 1176
rect -4032 1168 -4025 1176
rect -3982 1168 -3980 1176
rect -3975 1168 -3967 1176
rect -3960 1168 -3958 1176
rect -3330 1275 -3328 1283
rect -3323 1275 -3315 1283
rect -3308 1275 -3300 1283
rect -3295 1275 -3288 1283
rect -3922 1162 -3919 1171
rect -3915 1162 -3892 1171
rect -3888 1162 -3881 1171
rect -3849 1162 -3844 1171
rect -3839 1162 -3833 1171
rect -3722 1169 -3720 1177
rect -3715 1169 -3707 1177
rect -3700 1169 -3692 1177
rect -3687 1169 -3680 1177
rect -3637 1169 -3635 1177
rect -3630 1169 -3622 1177
rect -3615 1169 -3613 1177
rect -3407 1169 -3405 1177
rect -3400 1169 -3392 1177
rect -3385 1169 -3377 1177
rect -3372 1169 -3365 1177
rect -3322 1169 -3320 1177
rect -3315 1169 -3307 1177
rect -3300 1169 -3298 1177
rect -3262 1163 -3259 1172
rect -3255 1163 -3232 1172
rect -3228 1163 -3221 1172
rect -3189 1163 -3184 1172
rect -3179 1163 -3173 1172
rect -4658 1073 -4656 1081
rect -4651 1073 -4643 1081
rect -4636 1073 -4628 1081
rect -4623 1073 -4616 1081
rect -4573 1073 -4571 1081
rect -4566 1073 -4558 1081
rect -4551 1073 -4549 1081
rect -4277 1018 -4275 1026
rect -4270 1018 -4262 1026
rect -4255 1018 -4247 1026
rect -4242 1018 -4235 1026
rect -3990 1018 -3988 1026
rect -3983 1018 -3975 1026
rect -3968 1018 -3960 1026
rect -3955 1018 -3948 1026
rect -3644 1018 -3642 1026
rect -3637 1018 -3629 1026
rect -3622 1018 -3614 1026
rect -3609 1018 -3602 1026
rect -3362 1018 -3360 1026
rect -3355 1018 -3347 1026
rect -3340 1018 -3332 1026
rect -3327 1018 -3320 1026
rect -3035 1023 -3033 1031
rect -3028 1023 -3020 1031
rect -3013 1023 -3005 1031
rect -3000 1023 -2993 1031
rect -4658 966 -4656 974
rect -4651 966 -4643 974
rect -4636 966 -4628 974
rect -4623 966 -4616 974
rect -4573 966 -4571 974
rect -4566 966 -4558 974
rect -4551 966 -4549 974
rect -4358 943 -4356 951
rect -4351 943 -4343 951
rect -4336 943 -4328 951
rect -4323 943 -4316 951
rect -4191 940 -4189 948
rect -4184 940 -4176 948
rect -4169 940 -4161 948
rect -4156 940 -4149 948
rect -4071 943 -4069 951
rect -4064 943 -4056 951
rect -4049 943 -4041 951
rect -4036 943 -4029 951
rect -4658 866 -4656 874
rect -4651 866 -4643 874
rect -4636 866 -4628 874
rect -4623 866 -4616 874
rect -4573 866 -4571 874
rect -4566 866 -4558 874
rect -4551 866 -4549 874
rect -3904 940 -3902 948
rect -3897 940 -3889 948
rect -3882 940 -3874 948
rect -3869 940 -3862 948
rect -3725 943 -3723 951
rect -3718 943 -3710 951
rect -3703 943 -3695 951
rect -3690 943 -3683 951
rect -4277 858 -4275 866
rect -4270 858 -4262 866
rect -4255 858 -4247 866
rect -4242 858 -4235 866
rect -3558 940 -3556 948
rect -3551 940 -3543 948
rect -3536 940 -3528 948
rect -3523 940 -3516 948
rect -3443 943 -3441 951
rect -3436 943 -3428 951
rect -3421 943 -3413 951
rect -3408 943 -3401 951
rect -3990 858 -3988 866
rect -3983 858 -3975 866
rect -3968 858 -3960 866
rect -3955 858 -3948 866
rect -3116 948 -3114 956
rect -3109 948 -3101 956
rect -3094 948 -3086 956
rect -3081 948 -3074 956
rect -3276 940 -3274 948
rect -3269 940 -3261 948
rect -3254 940 -3246 948
rect -3241 940 -3234 948
rect -3644 858 -3642 866
rect -3637 858 -3629 866
rect -3622 858 -3614 866
rect -3609 858 -3602 866
rect -4659 751 -4657 759
rect -4652 751 -4644 759
rect -4637 751 -4629 759
rect -4624 751 -4617 759
rect -4574 751 -4572 759
rect -4567 751 -4559 759
rect -4552 751 -4550 759
rect -4354 752 -4352 760
rect -4347 752 -4339 760
rect -4332 752 -4324 760
rect -4319 752 -4312 760
rect -4269 752 -4267 760
rect -4262 752 -4254 760
rect -4247 752 -4245 760
rect -4067 752 -4065 760
rect -4060 752 -4052 760
rect -4045 752 -4037 760
rect -4032 752 -4025 760
rect -3982 752 -3980 760
rect -3975 752 -3967 760
rect -3960 752 -3958 760
rect -2949 945 -2947 953
rect -2942 945 -2934 953
rect -2927 945 -2919 953
rect -2914 945 -2907 953
rect -3362 858 -3360 866
rect -3355 858 -3347 866
rect -3340 858 -3332 866
rect -3327 858 -3320 866
rect -3035 863 -3033 871
rect -3028 863 -3020 871
rect -3013 863 -3005 871
rect -3000 863 -2993 871
rect -3922 746 -3919 755
rect -3915 746 -3892 755
rect -3888 746 -3881 755
rect -3849 746 -3844 755
rect -3839 746 -3833 755
rect -3721 752 -3719 760
rect -3714 752 -3706 760
rect -3699 752 -3691 760
rect -3686 752 -3679 760
rect -3636 752 -3634 760
rect -3629 752 -3621 760
rect -3614 752 -3612 760
rect -3439 752 -3437 760
rect -3432 752 -3424 760
rect -3417 752 -3409 760
rect -3404 752 -3397 760
rect -3354 752 -3352 760
rect -3347 752 -3339 760
rect -3332 752 -3330 760
rect -3112 757 -3110 765
rect -3105 757 -3097 765
rect -3090 757 -3082 765
rect -3077 757 -3070 765
rect -3027 757 -3025 765
rect -3020 757 -3012 765
rect -3005 757 -3003 765
rect -3294 746 -3291 755
rect -3287 746 -3264 755
rect -3260 746 -3253 755
rect -3221 746 -3216 755
rect -3211 746 -3205 755
rect -4659 651 -4657 659
rect -4652 651 -4644 659
rect -4637 651 -4629 659
rect -4624 651 -4617 659
rect -4574 651 -4572 659
rect -4567 651 -4559 659
rect -4552 651 -4550 659
rect -4277 560 -4275 568
rect -4270 560 -4262 568
rect -4255 560 -4247 568
rect -4242 560 -4235 568
rect -3978 560 -3976 568
rect -3971 560 -3963 568
rect -3956 560 -3948 568
rect -3943 560 -3936 568
rect -3663 560 -3661 568
rect -3656 560 -3648 568
rect -3641 560 -3633 568
rect -3628 560 -3621 568
rect -3334 566 -3332 574
rect -3327 566 -3319 574
rect -3312 566 -3304 574
rect -3299 566 -3292 574
rect -3019 566 -3017 574
rect -3012 566 -3004 574
rect -2997 566 -2989 574
rect -2984 566 -2977 574
rect -4659 544 -4657 552
rect -4652 544 -4644 552
rect -4637 544 -4629 552
rect -4624 544 -4617 552
rect -4574 544 -4572 552
rect -4567 544 -4559 552
rect -4552 544 -4550 552
rect -4358 485 -4356 493
rect -4351 485 -4343 493
rect -4336 485 -4328 493
rect -4323 485 -4316 493
rect -4659 444 -4657 452
rect -4652 444 -4644 452
rect -4637 444 -4629 452
rect -4624 444 -4617 452
rect -4574 444 -4572 452
rect -4567 444 -4559 452
rect -4552 444 -4550 452
rect -4191 482 -4189 490
rect -4184 482 -4176 490
rect -4169 482 -4161 490
rect -4156 482 -4149 490
rect -4059 485 -4057 493
rect -4052 485 -4044 493
rect -4037 485 -4029 493
rect -4024 485 -4017 493
rect -3892 482 -3890 490
rect -3885 482 -3877 490
rect -3870 482 -3862 490
rect -3857 482 -3850 490
rect -3744 485 -3742 493
rect -3737 485 -3729 493
rect -3722 485 -3714 493
rect -3709 485 -3702 493
rect -4277 400 -4275 408
rect -4270 400 -4262 408
rect -4255 400 -4247 408
rect -4242 400 -4235 408
rect -4659 341 -4657 349
rect -4652 341 -4644 349
rect -4637 341 -4629 349
rect -4624 341 -4617 349
rect -4574 341 -4572 349
rect -4567 341 -4559 349
rect -4552 341 -4550 349
rect -3415 491 -3413 499
rect -3408 491 -3400 499
rect -3393 491 -3385 499
rect -3380 491 -3373 499
rect -3577 482 -3575 490
rect -3570 482 -3562 490
rect -3555 482 -3547 490
rect -3542 482 -3535 490
rect -3978 400 -3976 408
rect -3971 400 -3963 408
rect -3956 400 -3948 408
rect -3943 400 -3936 408
rect -3248 488 -3246 496
rect -3241 488 -3233 496
rect -3226 488 -3218 496
rect -3213 488 -3206 496
rect -3100 491 -3098 499
rect -3093 491 -3085 499
rect -3078 491 -3070 499
rect -3065 491 -3058 499
rect -3663 400 -3661 408
rect -3656 400 -3648 408
rect -3641 400 -3633 408
rect -3628 400 -3621 408
rect -2933 488 -2931 496
rect -2926 488 -2918 496
rect -2911 488 -2903 496
rect -2898 488 -2891 496
rect -3334 406 -3332 414
rect -3327 406 -3319 414
rect -3312 406 -3304 414
rect -3299 406 -3292 414
rect -3019 406 -3017 414
rect -3012 406 -3004 414
rect -2997 406 -2989 414
rect -2984 406 -2977 414
rect -4354 294 -4352 302
rect -4347 294 -4339 302
rect -4332 294 -4324 302
rect -4319 294 -4312 302
rect -4269 294 -4267 302
rect -4262 294 -4254 302
rect -4247 294 -4245 302
rect -4055 294 -4053 302
rect -4048 294 -4040 302
rect -4033 294 -4025 302
rect -4020 294 -4013 302
rect -3970 294 -3968 302
rect -3963 294 -3955 302
rect -3948 294 -3946 302
rect -3740 294 -3738 302
rect -3733 294 -3725 302
rect -3718 294 -3710 302
rect -3705 294 -3698 302
rect -3655 294 -3653 302
rect -3648 294 -3640 302
rect -3633 294 -3631 302
rect -3411 300 -3409 308
rect -3404 300 -3396 308
rect -3389 300 -3381 308
rect -3376 300 -3369 308
rect -3326 300 -3324 308
rect -3319 300 -3311 308
rect -3304 300 -3302 308
rect -3096 300 -3094 308
rect -3089 300 -3081 308
rect -3074 300 -3066 308
rect -3061 300 -3054 308
rect -3011 300 -3009 308
rect -3004 300 -2996 308
rect -2989 300 -2987 308
rect -3595 268 -3592 277
rect -3588 268 -3565 277
rect -3561 268 -3554 277
rect -3522 268 -3517 277
rect -3512 268 -3506 277
rect -4659 241 -4657 249
rect -4652 241 -4644 249
rect -4637 241 -4629 249
rect -4624 241 -4617 249
rect -4574 241 -4572 249
rect -4567 241 -4559 249
rect -4552 241 -4550 249
rect -2951 274 -2948 283
rect -2944 274 -2921 283
rect -2917 274 -2910 283
rect -2878 274 -2873 283
rect -2868 274 -2862 283
rect -4277 186 -4275 194
rect -4270 186 -4262 194
rect -4255 186 -4247 194
rect -4242 186 -4235 194
rect -4659 134 -4657 142
rect -4652 134 -4644 142
rect -4637 134 -4629 142
rect -4624 134 -4617 142
rect -4574 134 -4572 142
rect -4567 134 -4559 142
rect -4552 134 -4550 142
rect -4358 111 -4356 119
rect -4351 111 -4343 119
rect -4336 111 -4328 119
rect -4323 111 -4316 119
rect -3946 153 -3944 161
rect -3939 153 -3931 161
rect -3924 153 -3916 161
rect -3911 153 -3904 161
rect -3631 153 -3629 161
rect -3624 153 -3616 161
rect -3609 153 -3601 161
rect -3596 153 -3589 161
rect -4191 108 -4189 116
rect -4184 108 -4176 116
rect -4169 108 -4161 116
rect -4156 108 -4149 116
rect -4659 34 -4657 42
rect -4652 34 -4644 42
rect -4637 34 -4629 42
rect -4624 34 -4617 42
rect -4574 34 -4572 42
rect -4567 34 -4559 42
rect -4552 34 -4550 42
rect -4027 78 -4025 86
rect -4020 78 -4012 86
rect -4005 78 -3997 86
rect -3992 78 -3985 86
rect -4277 26 -4275 34
rect -4270 26 -4262 34
rect -4255 26 -4247 34
rect -4242 26 -4235 34
rect -3860 75 -3858 83
rect -3853 75 -3845 83
rect -3838 75 -3830 83
rect -3825 75 -3818 83
rect -3712 78 -3710 86
rect -3705 78 -3697 86
rect -3690 78 -3682 86
rect -3677 78 -3670 86
rect -3545 75 -3543 83
rect -3538 75 -3530 83
rect -3523 75 -3515 83
rect -3510 75 -3503 83
rect -3946 -7 -3944 1
rect -3939 -7 -3931 1
rect -3924 -7 -3916 1
rect -3911 -7 -3904 1
rect -4354 -80 -4352 -72
rect -4347 -80 -4339 -72
rect -4332 -80 -4324 -72
rect -4319 -80 -4312 -72
rect -4269 -80 -4267 -72
rect -4262 -80 -4254 -72
rect -4247 -80 -4245 -72
rect -3631 -7 -3629 1
rect -3624 -7 -3616 1
rect -3609 -7 -3601 1
rect -3596 -7 -3589 1
rect -4023 -113 -4021 -105
rect -4016 -113 -4008 -105
rect -4001 -113 -3993 -105
rect -3988 -113 -3981 -105
rect -3938 -113 -3936 -105
rect -3931 -113 -3923 -105
rect -3916 -113 -3914 -105
rect -3708 -113 -3706 -105
rect -3701 -113 -3693 -105
rect -3686 -113 -3678 -105
rect -3673 -113 -3666 -105
rect -3623 -113 -3621 -105
rect -3616 -113 -3608 -105
rect -3601 -113 -3599 -105
rect -3563 -139 -3560 -130
rect -3556 -139 -3533 -130
rect -3529 -139 -3522 -130
rect -3490 -139 -3485 -130
rect -3480 -139 -3474 -130
rect -4277 -190 -4275 -182
rect -4270 -190 -4262 -182
rect -4255 -190 -4247 -182
rect -4242 -190 -4235 -182
rect -4358 -265 -4356 -257
rect -4351 -265 -4343 -257
rect -4336 -265 -4328 -257
rect -4323 -265 -4316 -257
rect -4191 -268 -4189 -260
rect -4184 -268 -4176 -260
rect -4169 -268 -4161 -260
rect -4156 -268 -4149 -260
rect -4277 -350 -4275 -342
rect -4270 -350 -4262 -342
rect -4255 -350 -4247 -342
rect -4242 -350 -4235 -342
rect -4354 -456 -4352 -448
rect -4347 -456 -4339 -448
rect -4332 -456 -4324 -448
rect -4319 -456 -4312 -448
rect -4269 -456 -4267 -448
rect -4262 -456 -4254 -448
rect -4247 -456 -4245 -448
<< ndcontact >>
rect -4646 1606 -4639 1612
rect -4622 1606 -4615 1612
rect -4573 1606 -4565 1612
rect -4555 1606 -4546 1612
rect -4670 1534 -4662 1543
rect -4616 1534 -4608 1543
rect -4587 1534 -4579 1543
rect -4558 1534 -4551 1543
rect -4646 1506 -4639 1512
rect -4619 1506 -4611 1512
rect -4573 1506 -4565 1512
rect -4555 1506 -4546 1512
rect -4265 1457 -4258 1464
rect -4244 1457 -4237 1464
rect -3978 1457 -3971 1464
rect -3957 1457 -3950 1464
rect -3633 1458 -3626 1465
rect -3612 1458 -3605 1465
rect -3318 1458 -3311 1465
rect -3297 1458 -3290 1465
rect -4670 1434 -4662 1443
rect -4616 1434 -4608 1443
rect -4587 1434 -4579 1443
rect -4558 1434 -4551 1443
rect -4646 1399 -4639 1405
rect -4573 1399 -4565 1405
rect -4555 1399 -4546 1405
rect -4346 1382 -4339 1389
rect -4325 1382 -4318 1389
rect -4289 1385 -4281 1394
rect -4235 1385 -4227 1394
rect -4670 1327 -4662 1336
rect -4616 1327 -4608 1336
rect -4587 1327 -4579 1336
rect -4558 1327 -4551 1336
rect -4646 1299 -4639 1305
rect -4179 1379 -4172 1386
rect -4158 1379 -4151 1386
rect -4059 1382 -4052 1389
rect -4038 1382 -4031 1389
rect -4002 1385 -3994 1394
rect -3948 1385 -3940 1394
rect -4370 1310 -4362 1319
rect -4316 1310 -4308 1319
rect -4619 1299 -4612 1305
rect -4573 1299 -4565 1305
rect -4555 1299 -4546 1305
rect -4265 1297 -4258 1304
rect -3892 1379 -3885 1386
rect -3871 1379 -3864 1386
rect -3714 1383 -3707 1390
rect -3693 1383 -3686 1390
rect -3657 1386 -3649 1395
rect -3603 1386 -3595 1395
rect -4203 1307 -4195 1316
rect -4149 1307 -4141 1316
rect -4083 1310 -4075 1319
rect -4029 1310 -4021 1319
rect -4241 1297 -4234 1304
rect -4670 1227 -4662 1236
rect -4616 1227 -4608 1236
rect -4587 1227 -4579 1236
rect -4558 1227 -4551 1236
rect -4646 1196 -4639 1202
rect -4623 1196 -4616 1202
rect -4573 1196 -4565 1202
rect -4555 1196 -4546 1202
rect -4342 1191 -4335 1197
rect -4321 1191 -4314 1197
rect -3978 1297 -3971 1304
rect -3547 1380 -3540 1387
rect -3526 1380 -3519 1387
rect -3399 1383 -3392 1390
rect -3378 1383 -3371 1390
rect -3342 1386 -3334 1395
rect -3288 1386 -3280 1395
rect -3916 1307 -3908 1316
rect -3862 1307 -3854 1316
rect -3738 1311 -3730 1320
rect -3684 1311 -3676 1320
rect -3954 1297 -3947 1304
rect -4289 1225 -4281 1234
rect -4235 1225 -4227 1234
rect -4269 1191 -4261 1197
rect -4251 1191 -4242 1197
rect -4055 1191 -4048 1197
rect -4034 1191 -4027 1197
rect -3633 1298 -3626 1305
rect -3232 1380 -3225 1387
rect -3211 1380 -3204 1387
rect -3571 1308 -3563 1317
rect -3517 1308 -3509 1317
rect -3423 1311 -3415 1320
rect -3369 1311 -3361 1320
rect -3609 1298 -3602 1305
rect -4002 1225 -3994 1234
rect -3948 1225 -3940 1234
rect -3982 1191 -3974 1197
rect -3964 1191 -3955 1197
rect -4670 1124 -4662 1133
rect -4616 1124 -4608 1133
rect -4587 1124 -4579 1133
rect -4558 1124 -4551 1133
rect -3918 1186 -3912 1192
rect -3710 1192 -3703 1198
rect -3689 1192 -3682 1198
rect -3892 1186 -3886 1192
rect -3865 1186 -3859 1192
rect -3846 1186 -3840 1192
rect -3318 1298 -3311 1305
rect -3256 1308 -3248 1317
rect -3202 1308 -3194 1317
rect -3294 1298 -3287 1305
rect -3657 1226 -3649 1235
rect -3603 1226 -3595 1235
rect -3637 1192 -3629 1198
rect -3619 1192 -3610 1198
rect -3395 1192 -3388 1198
rect -3374 1192 -3367 1198
rect -3342 1226 -3334 1235
rect -3288 1226 -3280 1235
rect -3322 1192 -3314 1198
rect -3304 1192 -3295 1198
rect -4646 1096 -4639 1102
rect -4366 1119 -4358 1128
rect -4312 1119 -4304 1128
rect -4283 1119 -4275 1128
rect -4254 1119 -4247 1128
rect -4079 1119 -4071 1128
rect -4025 1119 -4017 1128
rect -3996 1119 -3988 1128
rect -3967 1119 -3960 1128
rect -3258 1187 -3252 1193
rect -3232 1187 -3226 1193
rect -3205 1187 -3199 1193
rect -3186 1187 -3180 1193
rect -3928 1120 -3923 1125
rect -3908 1120 -3902 1125
rect -3882 1120 -3877 1125
rect -3859 1120 -3853 1125
rect -3833 1120 -3828 1125
rect -3734 1120 -3726 1129
rect -3680 1120 -3672 1129
rect -3651 1120 -3643 1129
rect -3622 1120 -3615 1129
rect -3419 1120 -3411 1129
rect -3365 1120 -3357 1129
rect -3336 1120 -3328 1129
rect -3307 1120 -3300 1129
rect -3268 1121 -3263 1126
rect -3248 1121 -3242 1126
rect -3222 1121 -3217 1126
rect -3199 1121 -3193 1126
rect -3173 1121 -3168 1126
rect -4619 1096 -4612 1102
rect -4573 1096 -4565 1102
rect -4555 1096 -4546 1102
rect -4265 1041 -4258 1048
rect -4244 1041 -4237 1048
rect -3978 1041 -3971 1048
rect -3957 1041 -3950 1048
rect -3632 1041 -3625 1048
rect -3611 1041 -3604 1048
rect -3350 1041 -3343 1048
rect -3329 1041 -3322 1048
rect -3023 1046 -3016 1053
rect -3002 1046 -2995 1053
rect -4670 1024 -4662 1033
rect -4616 1024 -4608 1033
rect -4587 1024 -4579 1033
rect -4558 1024 -4551 1033
rect -4646 989 -4639 995
rect -4620 989 -4612 995
rect -4573 989 -4565 995
rect -4555 989 -4546 995
rect -4346 966 -4339 973
rect -4325 966 -4318 973
rect -4289 969 -4281 978
rect -4235 969 -4227 978
rect -4670 917 -4662 926
rect -4616 917 -4608 926
rect -4587 917 -4579 926
rect -4558 917 -4551 926
rect -4646 889 -4639 895
rect -4179 963 -4172 970
rect -4158 963 -4151 970
rect -4059 966 -4052 973
rect -4038 966 -4031 973
rect -4002 969 -3994 978
rect -3948 969 -3940 978
rect -4620 889 -4612 895
rect -4573 889 -4565 895
rect -4555 889 -4546 895
rect -4370 894 -4362 903
rect -4316 894 -4308 903
rect -4265 881 -4258 888
rect -3892 963 -3885 970
rect -3871 963 -3864 970
rect -3713 966 -3706 973
rect -3692 966 -3685 973
rect -3656 969 -3648 978
rect -3602 969 -3594 978
rect -4203 891 -4195 900
rect -4149 891 -4141 900
rect -4083 894 -4075 903
rect -4029 894 -4021 903
rect -4241 881 -4234 888
rect -4670 817 -4662 826
rect -4616 817 -4608 826
rect -4587 817 -4579 826
rect -4558 817 -4551 826
rect -4647 774 -4640 780
rect -4623 774 -4616 780
rect -4574 774 -4566 780
rect -4556 774 -4547 780
rect -4342 775 -4335 781
rect -4321 775 -4314 781
rect -3978 881 -3971 888
rect -3546 963 -3539 970
rect -3525 963 -3518 970
rect -3431 966 -3424 973
rect -3410 966 -3403 973
rect -3374 969 -3366 978
rect -3320 969 -3312 978
rect -3916 891 -3908 900
rect -3862 891 -3854 900
rect -3737 894 -3729 903
rect -3683 894 -3675 903
rect -3954 881 -3947 888
rect -4289 809 -4281 818
rect -4235 809 -4227 818
rect -4269 775 -4261 781
rect -4251 775 -4242 781
rect -4055 775 -4048 781
rect -4034 775 -4027 781
rect -3632 881 -3625 888
rect -3264 963 -3257 970
rect -3243 963 -3236 970
rect -3104 971 -3097 978
rect -3083 971 -3076 978
rect -3047 974 -3039 983
rect -2993 974 -2985 983
rect -3570 891 -3562 900
rect -3516 891 -3508 900
rect -3455 894 -3447 903
rect -3401 894 -3393 903
rect -3608 881 -3601 888
rect -4002 809 -3994 818
rect -3948 809 -3940 818
rect -3982 775 -3974 781
rect -3964 775 -3955 781
rect -3918 770 -3912 776
rect -3892 770 -3886 776
rect -3865 770 -3859 776
rect -3846 770 -3840 776
rect -3709 775 -3702 781
rect -3688 775 -3681 781
rect -3350 881 -3343 888
rect -2937 968 -2930 975
rect -2916 968 -2909 975
rect -3288 891 -3280 900
rect -3234 891 -3226 900
rect -3128 899 -3120 908
rect -3074 899 -3066 908
rect -3326 881 -3319 888
rect -3656 809 -3648 818
rect -3602 809 -3594 818
rect -3636 775 -3628 781
rect -3618 775 -3609 781
rect -3427 775 -3420 781
rect -3406 775 -3399 781
rect -3023 886 -3016 893
rect -2961 896 -2953 905
rect -2907 896 -2899 905
rect -2999 886 -2992 893
rect -3374 809 -3366 818
rect -3320 809 -3312 818
rect -3354 775 -3346 781
rect -3336 775 -3327 781
rect -3100 780 -3093 786
rect -3079 780 -3072 786
rect -3047 814 -3039 823
rect -2993 814 -2985 823
rect -3027 780 -3019 786
rect -3009 780 -3000 786
rect -4671 702 -4663 711
rect -4617 702 -4609 711
rect -4588 702 -4580 711
rect -4559 702 -4552 711
rect -4366 703 -4358 712
rect -4312 703 -4304 712
rect -4283 703 -4275 712
rect -4254 703 -4247 712
rect -4079 703 -4071 712
rect -4025 703 -4017 712
rect -3996 703 -3988 712
rect -3967 703 -3960 712
rect -3290 770 -3284 776
rect -3264 770 -3258 776
rect -3237 770 -3231 776
rect -3218 770 -3212 776
rect -3928 704 -3923 709
rect -3908 704 -3902 709
rect -3882 704 -3877 709
rect -3859 704 -3853 709
rect -3833 704 -3828 709
rect -4647 674 -4640 680
rect -4622 674 -4614 680
rect -4574 674 -4566 680
rect -4556 674 -4547 680
rect -3733 703 -3725 712
rect -3679 703 -3671 712
rect -3650 703 -3642 712
rect -3621 703 -3614 712
rect -3451 703 -3443 712
rect -3397 703 -3389 712
rect -3368 703 -3360 712
rect -3339 703 -3332 712
rect -3300 704 -3295 709
rect -3280 704 -3274 709
rect -3254 704 -3249 709
rect -3231 704 -3225 709
rect -3205 704 -3200 709
rect -3124 708 -3116 717
rect -3070 708 -3062 717
rect -3041 708 -3033 717
rect -3012 708 -3005 717
rect -4671 602 -4663 611
rect -4617 602 -4609 611
rect -4588 602 -4580 611
rect -4559 602 -4552 611
rect -4647 567 -4640 573
rect -4265 583 -4258 590
rect -4244 583 -4237 590
rect -3966 583 -3959 590
rect -3945 583 -3938 590
rect -3651 583 -3644 590
rect -3630 583 -3623 590
rect -3322 589 -3315 596
rect -3301 589 -3294 596
rect -3007 589 -3000 596
rect -2986 589 -2979 596
rect -4622 567 -4615 573
rect -4574 567 -4566 573
rect -4556 567 -4547 573
rect -4671 495 -4663 504
rect -4617 495 -4609 504
rect -4588 495 -4580 504
rect -4559 495 -4552 504
rect -4647 467 -4640 473
rect -4346 508 -4339 515
rect -4322 508 -4315 515
rect -4289 511 -4281 520
rect -4235 511 -4227 520
rect -4622 467 -4615 473
rect -4574 467 -4566 473
rect -4556 467 -4547 473
rect -4179 505 -4172 512
rect -4158 505 -4151 512
rect -4047 508 -4040 515
rect -4026 508 -4019 515
rect -3990 511 -3982 520
rect -3936 511 -3928 520
rect -4370 436 -4362 445
rect -4316 436 -4308 445
rect -4671 395 -4663 404
rect -4617 395 -4609 404
rect -4588 395 -4580 404
rect -4559 395 -4552 404
rect -4265 423 -4258 430
rect -3880 505 -3873 512
rect -3859 505 -3852 512
rect -3732 508 -3725 515
rect -3711 508 -3704 515
rect -3675 511 -3667 520
rect -3621 511 -3613 520
rect -4203 433 -4195 442
rect -4149 433 -4141 442
rect -4071 436 -4063 445
rect -4017 436 -4009 445
rect -4241 423 -4234 430
rect -4647 364 -4640 370
rect -4624 364 -4617 370
rect -4574 364 -4566 370
rect -4556 364 -4547 370
rect -4342 317 -4335 323
rect -4321 317 -4314 323
rect -3966 423 -3959 430
rect -3565 505 -3558 512
rect -3544 505 -3537 512
rect -3403 514 -3396 521
rect -3382 514 -3375 521
rect -3346 517 -3338 526
rect -3292 517 -3284 526
rect -3904 433 -3896 442
rect -3850 433 -3842 442
rect -3756 436 -3748 445
rect -3702 436 -3694 445
rect -3942 423 -3935 430
rect -4289 351 -4281 360
rect -4235 351 -4227 360
rect -4269 317 -4261 323
rect -4251 317 -4242 323
rect -4043 317 -4036 323
rect -4022 317 -4015 323
rect -3651 423 -3644 430
rect -3236 511 -3229 518
rect -3215 511 -3208 518
rect -3088 514 -3081 521
rect -3067 514 -3060 521
rect -3031 517 -3023 526
rect -2977 517 -2969 526
rect -3427 442 -3419 451
rect -3373 442 -3365 451
rect -3589 433 -3581 442
rect -3535 433 -3527 442
rect -3627 423 -3620 430
rect -3990 351 -3982 360
rect -3936 351 -3928 360
rect -3970 317 -3962 323
rect -3952 317 -3943 323
rect -3728 317 -3721 323
rect -3707 317 -3700 323
rect -3322 429 -3315 436
rect -2921 511 -2914 518
rect -2900 511 -2893 518
rect -3260 439 -3252 448
rect -3206 439 -3198 448
rect -3112 442 -3104 451
rect -3058 442 -3050 451
rect -3298 429 -3291 436
rect -3675 351 -3667 360
rect -3621 351 -3613 360
rect -3399 323 -3392 329
rect -3378 323 -3371 329
rect -3655 317 -3647 323
rect -3637 317 -3628 323
rect -3007 429 -3000 436
rect -2945 439 -2937 448
rect -2891 439 -2883 448
rect -2983 429 -2976 436
rect -3346 357 -3338 366
rect -3292 357 -3284 366
rect -3326 323 -3318 329
rect -3308 323 -3299 329
rect -3084 323 -3077 329
rect -3063 323 -3056 329
rect -3031 357 -3023 366
rect -2977 357 -2969 366
rect -3011 323 -3003 329
rect -2993 323 -2984 329
rect -4671 292 -4663 301
rect -4617 292 -4609 301
rect -4588 292 -4580 301
rect -4559 292 -4552 301
rect -4647 264 -4640 270
rect -4622 264 -4615 270
rect -4574 264 -4566 270
rect -4556 264 -4547 270
rect -3591 292 -3585 298
rect -3565 292 -3559 298
rect -3538 292 -3532 298
rect -3519 292 -3513 298
rect -4366 245 -4358 254
rect -4312 245 -4304 254
rect -4283 245 -4275 254
rect -4254 245 -4247 254
rect -4067 245 -4059 254
rect -4013 245 -4005 254
rect -3984 245 -3976 254
rect -3955 245 -3948 254
rect -3752 245 -3744 254
rect -3698 245 -3690 254
rect -3669 245 -3661 254
rect -3640 245 -3633 254
rect -4265 209 -4258 216
rect -4244 209 -4237 216
rect -2947 298 -2941 304
rect -2921 298 -2915 304
rect -2894 298 -2888 304
rect -2875 298 -2869 304
rect -3423 251 -3415 260
rect -3369 251 -3361 260
rect -3340 251 -3332 260
rect -3311 251 -3304 260
rect -3108 251 -3100 260
rect -3054 251 -3046 260
rect -3025 251 -3017 260
rect -2996 251 -2989 260
rect -3601 226 -3596 231
rect -3581 226 -3575 231
rect -3555 226 -3550 231
rect -3532 226 -3526 231
rect -3506 226 -3501 231
rect -2957 232 -2952 237
rect -2937 232 -2931 237
rect -2911 232 -2906 237
rect -2888 232 -2882 237
rect -2862 232 -2857 237
rect -4671 192 -4663 201
rect -4617 192 -4609 201
rect -4588 192 -4580 201
rect -4559 192 -4552 201
rect -4647 157 -4640 163
rect -4622 157 -4615 163
rect -4574 157 -4566 163
rect -4556 157 -4547 163
rect -4346 134 -4339 141
rect -3934 176 -3927 183
rect -3913 176 -3906 183
rect -3619 176 -3612 183
rect -3598 176 -3591 183
rect -4321 134 -4314 141
rect -4289 137 -4281 146
rect -4235 137 -4227 146
rect -4671 85 -4663 94
rect -4617 85 -4609 94
rect -4588 85 -4580 94
rect -4559 85 -4552 94
rect -4647 57 -4640 63
rect -4179 131 -4172 138
rect -4158 131 -4151 138
rect -4623 57 -4616 63
rect -4574 57 -4566 63
rect -4556 57 -4547 63
rect -4370 62 -4362 71
rect -4316 62 -4308 71
rect -4265 49 -4258 56
rect -4015 101 -4008 108
rect -3994 101 -3987 108
rect -3958 104 -3950 113
rect -3904 104 -3896 113
rect -4203 59 -4195 68
rect -4149 59 -4141 68
rect -4241 49 -4234 56
rect -4671 -15 -4663 -6
rect -4617 -15 -4609 -6
rect -4588 -15 -4580 -6
rect -4559 -15 -4552 -6
rect -4342 -57 -4335 -51
rect -4321 -57 -4314 -51
rect -3848 98 -3841 105
rect -3827 98 -3820 105
rect -3700 101 -3693 108
rect -3679 101 -3672 108
rect -3643 104 -3635 113
rect -3589 104 -3581 113
rect -4039 29 -4031 38
rect -3985 29 -3977 38
rect -4289 -23 -4281 -14
rect -4235 -23 -4227 -14
rect -3934 16 -3927 23
rect -3533 98 -3526 105
rect -3512 98 -3505 105
rect -3872 26 -3864 35
rect -3818 26 -3810 35
rect -3724 29 -3716 38
rect -3670 29 -3662 38
rect -3910 16 -3903 23
rect -4269 -57 -4261 -51
rect -4251 -57 -4242 -51
rect -4011 -90 -4004 -84
rect -3990 -90 -3983 -84
rect -3619 16 -3612 23
rect -3557 26 -3549 35
rect -3503 26 -3495 35
rect -3595 16 -3588 23
rect -3958 -56 -3950 -47
rect -3904 -56 -3896 -47
rect -3938 -90 -3930 -84
rect -3920 -90 -3911 -84
rect -3696 -90 -3689 -84
rect -3675 -90 -3668 -84
rect -3643 -56 -3635 -47
rect -3589 -56 -3581 -47
rect -3623 -90 -3615 -84
rect -3605 -90 -3596 -84
rect -4366 -129 -4358 -120
rect -4312 -129 -4304 -120
rect -4283 -129 -4275 -120
rect -4254 -129 -4247 -120
rect -3559 -115 -3553 -109
rect -3533 -115 -3527 -109
rect -3506 -115 -3500 -109
rect -3487 -115 -3481 -109
rect -4265 -167 -4258 -160
rect -4244 -167 -4237 -160
rect -4035 -162 -4027 -153
rect -3981 -162 -3973 -153
rect -3952 -162 -3944 -153
rect -3923 -162 -3916 -153
rect -3720 -162 -3712 -153
rect -3666 -162 -3658 -153
rect -3637 -162 -3629 -153
rect -3608 -162 -3601 -153
rect -4346 -242 -4339 -235
rect -3569 -181 -3564 -176
rect -3549 -181 -3543 -176
rect -3523 -181 -3518 -176
rect -3500 -181 -3494 -176
rect -3474 -181 -3469 -176
rect -4321 -242 -4314 -235
rect -4289 -239 -4281 -230
rect -4235 -239 -4227 -230
rect -4179 -245 -4172 -238
rect -4158 -245 -4151 -238
rect -4370 -314 -4362 -305
rect -4316 -314 -4308 -305
rect -4265 -327 -4258 -320
rect -4203 -317 -4195 -308
rect -4149 -317 -4141 -308
rect -4241 -327 -4234 -320
rect -4342 -433 -4335 -427
rect -4321 -433 -4314 -427
rect -4289 -399 -4281 -390
rect -4235 -399 -4227 -390
rect -4269 -433 -4261 -427
rect -4251 -433 -4242 -427
rect -4366 -505 -4358 -496
rect -4312 -505 -4304 -496
rect -4283 -505 -4275 -496
rect -4254 -505 -4247 -496
<< pdcontact >>
rect -4665 1583 -4658 1591
rect -4643 1583 -4636 1591
rect -4616 1583 -4609 1591
rect -4580 1583 -4573 1591
rect -4558 1583 -4551 1591
rect -4665 1483 -4658 1491
rect -4643 1483 -4636 1491
rect -4616 1483 -4609 1491
rect -4580 1483 -4573 1491
rect -4558 1483 -4551 1491
rect -4284 1434 -4277 1442
rect -4262 1434 -4255 1442
rect -4235 1434 -4228 1442
rect -3997 1434 -3990 1442
rect -3975 1434 -3968 1442
rect -3948 1434 -3941 1442
rect -3652 1435 -3645 1443
rect -3630 1435 -3623 1443
rect -3603 1435 -3596 1443
rect -3337 1435 -3330 1443
rect -3315 1435 -3308 1443
rect -3288 1435 -3281 1443
rect -4665 1376 -4658 1384
rect -4643 1376 -4636 1384
rect -4616 1376 -4609 1384
rect -4580 1376 -4573 1384
rect -4558 1376 -4551 1384
rect -4365 1359 -4358 1367
rect -4343 1359 -4336 1367
rect -4316 1359 -4309 1367
rect -4198 1356 -4191 1364
rect -4176 1356 -4169 1364
rect -4149 1356 -4142 1364
rect -4078 1359 -4071 1367
rect -4056 1359 -4049 1367
rect -4029 1359 -4022 1367
rect -4665 1276 -4658 1284
rect -4643 1276 -4636 1284
rect -4616 1276 -4609 1284
rect -4580 1276 -4573 1284
rect -4558 1276 -4551 1284
rect -3911 1356 -3904 1364
rect -3889 1356 -3882 1364
rect -3862 1356 -3855 1364
rect -3733 1360 -3726 1368
rect -3711 1360 -3704 1368
rect -3684 1360 -3677 1368
rect -4284 1274 -4277 1282
rect -4262 1274 -4255 1282
rect -4235 1274 -4228 1282
rect -3566 1357 -3559 1365
rect -3544 1357 -3537 1365
rect -3517 1357 -3510 1365
rect -3418 1360 -3411 1368
rect -3396 1360 -3389 1368
rect -3369 1360 -3362 1368
rect -3997 1274 -3990 1282
rect -3975 1274 -3968 1282
rect -3948 1274 -3941 1282
rect -3251 1357 -3244 1365
rect -3229 1357 -3222 1365
rect -3202 1357 -3195 1365
rect -3652 1275 -3645 1283
rect -3630 1275 -3623 1283
rect -3603 1275 -3596 1283
rect -4665 1173 -4658 1181
rect -4643 1173 -4636 1181
rect -4616 1173 -4609 1181
rect -4580 1173 -4573 1181
rect -4558 1173 -4551 1181
rect -4361 1168 -4354 1176
rect -4339 1168 -4332 1176
rect -4312 1168 -4305 1176
rect -4276 1168 -4269 1176
rect -4254 1168 -4247 1176
rect -4074 1168 -4067 1176
rect -4052 1168 -4045 1176
rect -4025 1168 -4018 1176
rect -3989 1168 -3982 1176
rect -3967 1168 -3960 1176
rect -3337 1275 -3330 1283
rect -3315 1275 -3308 1283
rect -3288 1275 -3281 1283
rect -3927 1162 -3922 1171
rect -3881 1162 -3876 1171
rect -3854 1162 -3849 1171
rect -3833 1162 -3828 1171
rect -3729 1169 -3722 1177
rect -3707 1169 -3700 1177
rect -3680 1169 -3673 1177
rect -3644 1169 -3637 1177
rect -3622 1169 -3615 1177
rect -3414 1169 -3407 1177
rect -3392 1169 -3385 1177
rect -3365 1169 -3358 1177
rect -3329 1169 -3322 1177
rect -3307 1169 -3300 1177
rect -3267 1163 -3262 1172
rect -3221 1163 -3216 1172
rect -3194 1163 -3189 1172
rect -3173 1163 -3168 1172
rect -3922 1102 -3916 1108
rect -3891 1102 -3885 1108
rect -3869 1102 -3863 1108
rect -3850 1102 -3844 1108
rect -3262 1103 -3256 1109
rect -3231 1103 -3225 1109
rect -3209 1103 -3203 1109
rect -3190 1103 -3184 1109
rect -4665 1073 -4658 1081
rect -4643 1073 -4636 1081
rect -4616 1073 -4609 1081
rect -4580 1073 -4573 1081
rect -4558 1073 -4551 1081
rect -4284 1018 -4277 1026
rect -4262 1018 -4255 1026
rect -4235 1018 -4228 1026
rect -3997 1018 -3990 1026
rect -3975 1018 -3968 1026
rect -3948 1018 -3941 1026
rect -3651 1018 -3644 1026
rect -3629 1018 -3622 1026
rect -3602 1018 -3595 1026
rect -3369 1018 -3362 1026
rect -3347 1018 -3340 1026
rect -3320 1018 -3313 1026
rect -3042 1023 -3035 1031
rect -3020 1023 -3013 1031
rect -2993 1023 -2986 1031
rect -4665 966 -4658 974
rect -4643 966 -4636 974
rect -4616 966 -4609 974
rect -4580 966 -4573 974
rect -4558 966 -4551 974
rect -4365 943 -4358 951
rect -4343 943 -4336 951
rect -4316 943 -4309 951
rect -4198 940 -4191 948
rect -4176 940 -4169 948
rect -4149 940 -4142 948
rect -4078 943 -4071 951
rect -4056 943 -4049 951
rect -4029 943 -4022 951
rect -4665 866 -4658 874
rect -4643 866 -4636 874
rect -4616 866 -4609 874
rect -4580 866 -4573 874
rect -4558 866 -4551 874
rect -3911 940 -3904 948
rect -3889 940 -3882 948
rect -3862 940 -3855 948
rect -3732 943 -3725 951
rect -3710 943 -3703 951
rect -3683 943 -3676 951
rect -4284 858 -4277 866
rect -4262 858 -4255 866
rect -4235 858 -4228 866
rect -3565 940 -3558 948
rect -3543 940 -3536 948
rect -3516 940 -3509 948
rect -3450 943 -3443 951
rect -3428 943 -3421 951
rect -3401 943 -3394 951
rect -3997 858 -3990 866
rect -3975 858 -3968 866
rect -3948 858 -3941 866
rect -3123 948 -3116 956
rect -3101 948 -3094 956
rect -3074 948 -3067 956
rect -3283 940 -3276 948
rect -3261 940 -3254 948
rect -3234 940 -3227 948
rect -3651 858 -3644 866
rect -3629 858 -3622 866
rect -3602 858 -3595 866
rect -4666 751 -4659 759
rect -4644 751 -4637 759
rect -4617 751 -4610 759
rect -4581 751 -4574 759
rect -4559 751 -4552 759
rect -4361 752 -4354 760
rect -4339 752 -4332 760
rect -4312 752 -4305 760
rect -4276 752 -4269 760
rect -4254 752 -4247 760
rect -4074 752 -4067 760
rect -4052 752 -4045 760
rect -4025 752 -4018 760
rect -3989 752 -3982 760
rect -3967 752 -3960 760
rect -2956 945 -2949 953
rect -2934 945 -2927 953
rect -2907 945 -2900 953
rect -3369 858 -3362 866
rect -3347 858 -3340 866
rect -3320 858 -3313 866
rect -3042 863 -3035 871
rect -3020 863 -3013 871
rect -2993 863 -2986 871
rect -3927 746 -3922 755
rect -3881 746 -3876 755
rect -3854 746 -3849 755
rect -3833 746 -3828 755
rect -3728 752 -3721 760
rect -3706 752 -3699 760
rect -3679 752 -3672 760
rect -3643 752 -3636 760
rect -3621 752 -3614 760
rect -3446 752 -3439 760
rect -3424 752 -3417 760
rect -3397 752 -3390 760
rect -3361 752 -3354 760
rect -3339 752 -3332 760
rect -3119 757 -3112 765
rect -3097 757 -3090 765
rect -3070 757 -3063 765
rect -3034 757 -3027 765
rect -3012 757 -3005 765
rect -3299 746 -3294 755
rect -3253 746 -3248 755
rect -3226 746 -3221 755
rect -3205 746 -3200 755
rect -3922 686 -3916 692
rect -3891 686 -3885 692
rect -3869 686 -3863 692
rect -3850 686 -3844 692
rect -3294 686 -3288 692
rect -3263 686 -3257 692
rect -3241 686 -3235 692
rect -3222 686 -3216 692
rect -4666 651 -4659 659
rect -4644 651 -4637 659
rect -4617 651 -4610 659
rect -4581 651 -4574 659
rect -4559 651 -4552 659
rect -4284 560 -4277 568
rect -4262 560 -4255 568
rect -4235 560 -4228 568
rect -3985 560 -3978 568
rect -3963 560 -3956 568
rect -3936 560 -3929 568
rect -3670 560 -3663 568
rect -3648 560 -3641 568
rect -3621 560 -3614 568
rect -3341 566 -3334 574
rect -3319 566 -3312 574
rect -3292 566 -3285 574
rect -3026 566 -3019 574
rect -3004 566 -2997 574
rect -2977 566 -2970 574
rect -4666 544 -4659 552
rect -4644 544 -4637 552
rect -4617 544 -4610 552
rect -4581 544 -4574 552
rect -4559 544 -4552 552
rect -4365 485 -4358 493
rect -4343 485 -4336 493
rect -4316 485 -4309 493
rect -4666 444 -4659 452
rect -4644 444 -4637 452
rect -4617 444 -4610 452
rect -4581 444 -4574 452
rect -4559 444 -4552 452
rect -4198 482 -4191 490
rect -4176 482 -4169 490
rect -4149 482 -4142 490
rect -4066 485 -4059 493
rect -4044 485 -4037 493
rect -4017 485 -4010 493
rect -3899 482 -3892 490
rect -3877 482 -3870 490
rect -3850 482 -3843 490
rect -3751 485 -3744 493
rect -3729 485 -3722 493
rect -3702 485 -3695 493
rect -4284 400 -4277 408
rect -4262 400 -4255 408
rect -4235 400 -4228 408
rect -4666 341 -4659 349
rect -4644 341 -4637 349
rect -4617 341 -4610 349
rect -4581 341 -4574 349
rect -4559 341 -4552 349
rect -3422 491 -3415 499
rect -3400 491 -3393 499
rect -3373 491 -3366 499
rect -3584 482 -3577 490
rect -3562 482 -3555 490
rect -3535 482 -3528 490
rect -3985 400 -3978 408
rect -3963 400 -3956 408
rect -3936 400 -3929 408
rect -3255 488 -3248 496
rect -3233 488 -3226 496
rect -3206 488 -3199 496
rect -3107 491 -3100 499
rect -3085 491 -3078 499
rect -3058 491 -3051 499
rect -3670 400 -3663 408
rect -3648 400 -3641 408
rect -3621 400 -3614 408
rect -2940 488 -2933 496
rect -2918 488 -2911 496
rect -2891 488 -2884 496
rect -3341 406 -3334 414
rect -3319 406 -3312 414
rect -3292 406 -3285 414
rect -3026 406 -3019 414
rect -3004 406 -2997 414
rect -2977 406 -2970 414
rect -4361 294 -4354 302
rect -4339 294 -4332 302
rect -4312 294 -4305 302
rect -4276 294 -4269 302
rect -4254 294 -4247 302
rect -4062 294 -4055 302
rect -4040 294 -4033 302
rect -4013 294 -4006 302
rect -3977 294 -3970 302
rect -3955 294 -3948 302
rect -3747 294 -3740 302
rect -3725 294 -3718 302
rect -3698 294 -3691 302
rect -3662 294 -3655 302
rect -3640 294 -3633 302
rect -3418 300 -3411 308
rect -3396 300 -3389 308
rect -3369 300 -3362 308
rect -3333 300 -3326 308
rect -3311 300 -3304 308
rect -3103 300 -3096 308
rect -3081 300 -3074 308
rect -3054 300 -3047 308
rect -3018 300 -3011 308
rect -2996 300 -2989 308
rect -3600 268 -3595 277
rect -3554 268 -3549 277
rect -3527 268 -3522 277
rect -3506 268 -3501 277
rect -4666 241 -4659 249
rect -4644 241 -4637 249
rect -4617 241 -4610 249
rect -4581 241 -4574 249
rect -4559 241 -4552 249
rect -2956 274 -2951 283
rect -2910 274 -2905 283
rect -2883 274 -2878 283
rect -2862 274 -2857 283
rect -3595 208 -3589 214
rect -3564 208 -3558 214
rect -3542 208 -3536 214
rect -3523 208 -3517 214
rect -2951 214 -2945 220
rect -2920 214 -2914 220
rect -2898 214 -2892 220
rect -2879 214 -2873 220
rect -4284 186 -4277 194
rect -4262 186 -4255 194
rect -4235 186 -4228 194
rect -4666 134 -4659 142
rect -4644 134 -4637 142
rect -4617 134 -4610 142
rect -4581 134 -4574 142
rect -4559 134 -4552 142
rect -4365 111 -4358 119
rect -4343 111 -4336 119
rect -4316 111 -4309 119
rect -3953 153 -3946 161
rect -3931 153 -3924 161
rect -3904 153 -3897 161
rect -3638 153 -3631 161
rect -3616 153 -3609 161
rect -3589 153 -3582 161
rect -4198 108 -4191 116
rect -4176 108 -4169 116
rect -4149 108 -4142 116
rect -4666 34 -4659 42
rect -4644 34 -4637 42
rect -4617 34 -4610 42
rect -4581 34 -4574 42
rect -4559 34 -4552 42
rect -4034 78 -4027 86
rect -4012 78 -4005 86
rect -3985 78 -3978 86
rect -4284 26 -4277 34
rect -4262 26 -4255 34
rect -4235 26 -4228 34
rect -3867 75 -3860 83
rect -3845 75 -3838 83
rect -3818 75 -3811 83
rect -3719 78 -3712 86
rect -3697 78 -3690 86
rect -3670 78 -3663 86
rect -3552 75 -3545 83
rect -3530 75 -3523 83
rect -3503 75 -3496 83
rect -3953 -7 -3946 1
rect -3931 -7 -3924 1
rect -3904 -7 -3897 1
rect -4361 -80 -4354 -72
rect -4339 -80 -4332 -72
rect -4312 -80 -4305 -72
rect -4276 -80 -4269 -72
rect -4254 -80 -4247 -72
rect -3638 -7 -3631 1
rect -3616 -7 -3609 1
rect -3589 -7 -3582 1
rect -4030 -113 -4023 -105
rect -4008 -113 -4001 -105
rect -3981 -113 -3974 -105
rect -3945 -113 -3938 -105
rect -3923 -113 -3916 -105
rect -3715 -113 -3708 -105
rect -3693 -113 -3686 -105
rect -3666 -113 -3659 -105
rect -3630 -113 -3623 -105
rect -3608 -113 -3601 -105
rect -3568 -139 -3563 -130
rect -3522 -139 -3517 -130
rect -3495 -139 -3490 -130
rect -3474 -139 -3469 -130
rect -4284 -190 -4277 -182
rect -4262 -190 -4255 -182
rect -4235 -190 -4228 -182
rect -3563 -199 -3557 -193
rect -3532 -199 -3526 -193
rect -3510 -199 -3504 -193
rect -3491 -199 -3485 -193
rect -4365 -265 -4358 -257
rect -4343 -265 -4336 -257
rect -4316 -265 -4309 -257
rect -4198 -268 -4191 -260
rect -4176 -268 -4169 -260
rect -4149 -268 -4142 -260
rect -4284 -350 -4277 -342
rect -4262 -350 -4255 -342
rect -4235 -350 -4228 -342
rect -4361 -456 -4354 -448
rect -4339 -456 -4332 -448
rect -4312 -456 -4305 -448
rect -4276 -456 -4269 -448
rect -4254 -456 -4247 -448
<< psubstratepcontact >>
rect -4658 1517 -4650 1525
rect -4622 1517 -4614 1525
rect -4579 1517 -4570 1525
rect -4560 1517 -4551 1525
rect -4658 1417 -4650 1425
rect -4622 1417 -4614 1425
rect -4579 1417 -4570 1425
rect -4560 1417 -4551 1425
rect -4277 1368 -4269 1376
rect -4658 1310 -4650 1318
rect -3990 1368 -3982 1376
rect -4622 1310 -4614 1318
rect -4579 1310 -4570 1318
rect -4560 1310 -4551 1318
rect -4358 1293 -4350 1301
rect -3645 1369 -3637 1377
rect -4191 1290 -4183 1298
rect -4658 1210 -4650 1218
rect -4622 1210 -4614 1218
rect -4579 1210 -4570 1218
rect -4560 1210 -4551 1218
rect -4071 1293 -4063 1301
rect -3330 1369 -3322 1377
rect -3904 1290 -3896 1298
rect -4277 1208 -4269 1216
rect -4249 1208 -4241 1216
rect -3726 1294 -3718 1302
rect -3559 1291 -3551 1299
rect -3990 1208 -3982 1216
rect -3962 1208 -3954 1216
rect -3411 1294 -3403 1302
rect -3244 1291 -3236 1299
rect -3645 1209 -3637 1217
rect -3617 1209 -3609 1217
rect -3330 1209 -3322 1217
rect -3302 1209 -3294 1217
rect -4658 1107 -4650 1115
rect -4622 1107 -4614 1115
rect -4579 1107 -4570 1115
rect -4560 1107 -4551 1115
rect -4354 1102 -4346 1110
rect -4317 1102 -4309 1110
rect -4275 1102 -4266 1110
rect -4256 1102 -4247 1110
rect -4067 1102 -4059 1110
rect -4031 1102 -4023 1110
rect -3988 1102 -3979 1110
rect -3969 1102 -3960 1110
rect -3722 1103 -3714 1111
rect -3685 1103 -3677 1111
rect -3643 1103 -3634 1111
rect -3624 1103 -3615 1111
rect -3407 1103 -3399 1111
rect -3371 1103 -3363 1111
rect -3328 1103 -3319 1111
rect -3309 1103 -3300 1111
rect -4658 1007 -4650 1015
rect -4622 1007 -4614 1015
rect -4579 1007 -4570 1015
rect -4560 1007 -4551 1015
rect -4277 952 -4269 960
rect -4658 900 -4650 908
rect -4622 900 -4614 908
rect -4579 900 -4570 908
rect -4560 900 -4551 908
rect -3990 952 -3982 960
rect -4358 877 -4350 885
rect -3644 952 -3636 960
rect -4191 874 -4183 882
rect -4658 800 -4650 808
rect -4622 800 -4614 808
rect -4579 800 -4570 808
rect -4560 800 -4551 808
rect -4071 877 -4063 885
rect -3362 952 -3354 960
rect -3904 874 -3896 882
rect -4277 792 -4269 800
rect -4249 792 -4241 800
rect -3725 877 -3717 885
rect -3035 957 -3027 965
rect -3558 874 -3550 882
rect -3990 792 -3982 800
rect -3962 792 -3954 800
rect -3443 877 -3435 885
rect -3276 874 -3268 882
rect -3644 792 -3636 800
rect -3616 792 -3608 800
rect -3116 882 -3108 890
rect -2949 879 -2941 887
rect -3362 792 -3354 800
rect -3334 792 -3326 800
rect -3035 797 -3027 805
rect -3007 797 -2999 805
rect -4659 685 -4651 693
rect -4623 685 -4615 693
rect -4580 685 -4571 693
rect -4561 685 -4552 693
rect -4354 686 -4346 694
rect -4317 686 -4309 694
rect -4275 686 -4266 694
rect -4256 686 -4247 694
rect -4067 686 -4059 694
rect -4031 686 -4023 694
rect -3988 686 -3979 694
rect -3969 686 -3960 694
rect -3721 686 -3713 694
rect -3684 686 -3676 694
rect -3642 686 -3633 694
rect -3623 686 -3614 694
rect -3439 686 -3431 694
rect -3403 686 -3395 694
rect -3360 686 -3351 694
rect -3341 686 -3332 694
rect -3112 691 -3104 699
rect -3074 691 -3066 699
rect -3033 691 -3024 699
rect -3014 691 -3005 699
rect -4659 585 -4651 593
rect -4623 585 -4615 593
rect -4580 585 -4571 593
rect -4561 585 -4552 593
rect -4659 478 -4651 486
rect -4277 494 -4269 502
rect -4623 478 -4615 486
rect -4580 478 -4571 486
rect -4561 478 -4552 486
rect -3978 494 -3970 502
rect -4358 419 -4350 427
rect -3663 494 -3655 502
rect -4191 416 -4183 424
rect -4659 378 -4651 386
rect -4623 378 -4615 386
rect -4580 378 -4571 386
rect -4561 378 -4552 386
rect -4059 419 -4051 427
rect -3334 500 -3326 508
rect -3892 416 -3884 424
rect -4277 334 -4269 342
rect -4249 334 -4241 342
rect -3744 419 -3736 427
rect -3019 500 -3011 508
rect -3577 416 -3569 424
rect -3978 334 -3970 342
rect -3950 334 -3942 342
rect -3415 425 -3407 433
rect -3248 422 -3240 430
rect -3663 334 -3655 342
rect -3635 334 -3627 342
rect -3100 425 -3092 433
rect -2933 422 -2925 430
rect -3334 340 -3326 348
rect -3306 340 -3298 348
rect -3019 340 -3011 348
rect -2991 340 -2983 348
rect -4659 275 -4651 283
rect -4623 275 -4615 283
rect -4580 275 -4571 283
rect -4561 275 -4552 283
rect -4354 228 -4346 236
rect -4326 228 -4318 236
rect -4275 228 -4266 236
rect -4256 228 -4247 236
rect -4055 228 -4047 236
rect -4018 228 -4010 236
rect -3976 228 -3967 236
rect -3957 228 -3948 236
rect -3740 228 -3732 236
rect -3703 228 -3695 236
rect -3661 228 -3652 236
rect -3642 228 -3633 236
rect -3411 234 -3403 242
rect -3374 234 -3366 242
rect -3332 234 -3323 242
rect -3313 234 -3304 242
rect -3096 234 -3088 242
rect -3060 234 -3052 242
rect -3017 234 -3008 242
rect -2998 234 -2989 242
rect -4659 175 -4651 183
rect -4623 175 -4615 183
rect -4580 175 -4571 183
rect -4561 175 -4552 183
rect -4277 120 -4269 128
rect -4659 68 -4651 76
rect -4623 68 -4615 76
rect -4580 68 -4571 76
rect -4561 68 -4552 76
rect -4358 45 -4350 53
rect -3946 87 -3938 95
rect -4191 42 -4183 50
rect -4659 -32 -4651 -24
rect -4623 -32 -4615 -24
rect -4580 -32 -4571 -24
rect -4561 -32 -4552 -24
rect -3631 87 -3623 95
rect -4027 12 -4019 20
rect -3860 9 -3852 17
rect -4277 -40 -4269 -32
rect -4249 -40 -4241 -32
rect -3712 12 -3704 20
rect -3545 9 -3537 17
rect -3946 -73 -3938 -65
rect -3918 -73 -3910 -65
rect -3631 -73 -3623 -65
rect -3603 -73 -3595 -65
rect -4354 -146 -4346 -138
rect -4326 -146 -4318 -138
rect -4275 -146 -4266 -138
rect -4256 -146 -4247 -138
rect -4023 -179 -4015 -171
rect -3986 -179 -3978 -171
rect -3944 -179 -3935 -171
rect -3925 -179 -3916 -171
rect -3708 -179 -3700 -171
rect -3672 -179 -3664 -171
rect -3629 -179 -3620 -171
rect -3610 -179 -3601 -171
rect -4277 -256 -4269 -248
rect -4358 -331 -4350 -323
rect -4191 -334 -4183 -326
rect -4277 -416 -4269 -408
rect -4249 -416 -4241 -408
rect -4354 -522 -4346 -514
rect -4326 -522 -4318 -514
rect -4275 -522 -4266 -514
rect -4256 -522 -4247 -514
<< polysilicon >>
rect -4656 1591 -4651 1599
rect -4628 1591 -4623 1599
rect -4571 1591 -4566 1599
rect -4656 1559 -4651 1583
rect -4702 1553 -4651 1559
rect -4656 1543 -4651 1553
rect -4628 1543 -4623 1583
rect -4571 1567 -4566 1583
rect -4608 1559 -4566 1567
rect -4571 1543 -4566 1559
rect -4656 1531 -4651 1534
rect -4656 1491 -4651 1499
rect -4628 1491 -4623 1534
rect -4571 1530 -4566 1534
rect -4571 1491 -4566 1499
rect -4656 1456 -4651 1483
rect -4693 1450 -4651 1456
rect -4656 1443 -4651 1450
rect -4628 1443 -4623 1483
rect -4571 1467 -4566 1483
rect -4608 1459 -4566 1467
rect -4571 1443 -4566 1459
rect -4275 1442 -4270 1450
rect -4247 1442 -4242 1450
rect -3988 1442 -3983 1450
rect -3960 1442 -3955 1450
rect -3643 1443 -3638 1451
rect -3615 1443 -3610 1451
rect -3328 1443 -3323 1451
rect -3300 1443 -3295 1451
rect -4656 1431 -4651 1434
rect -4656 1384 -4651 1392
rect -4628 1384 -4623 1434
rect -4571 1430 -4566 1434
rect -4275 1417 -4270 1434
rect -4356 1412 -4352 1417
rect -4281 1412 -4270 1417
rect -4571 1384 -4566 1392
rect -4656 1354 -4651 1376
rect -4684 1348 -4651 1354
rect -4656 1336 -4651 1348
rect -4628 1336 -4623 1376
rect -4571 1360 -4566 1376
rect -4356 1367 -4351 1412
rect -4275 1394 -4270 1412
rect -4247 1394 -4242 1434
rect -4227 1410 -4222 1418
rect -3988 1417 -3983 1434
rect -4275 1382 -4270 1385
rect -4328 1367 -4323 1375
rect -4608 1352 -4566 1360
rect -4571 1336 -4566 1352
rect -4356 1334 -4351 1359
rect -4375 1327 -4351 1334
rect -4656 1324 -4651 1327
rect -4656 1284 -4651 1292
rect -4628 1284 -4623 1327
rect -4571 1323 -4566 1327
rect -4356 1319 -4351 1327
rect -4328 1319 -4323 1359
rect -4247 1343 -4242 1385
rect -4189 1364 -4184 1410
rect -4069 1412 -4065 1417
rect -3994 1412 -3983 1417
rect -4161 1364 -4156 1372
rect -4069 1367 -4064 1412
rect -3988 1394 -3983 1412
rect -3960 1394 -3955 1434
rect -3643 1418 -3638 1435
rect -3940 1410 -3935 1418
rect -3988 1382 -3983 1385
rect -4041 1367 -4036 1375
rect -4308 1335 -4242 1343
rect -4356 1307 -4351 1310
rect -4571 1284 -4566 1292
rect -4656 1254 -4651 1276
rect -4675 1248 -4651 1254
rect -4656 1236 -4651 1248
rect -4628 1236 -4623 1276
rect -4571 1260 -4566 1276
rect -4608 1252 -4566 1260
rect -4571 1236 -4566 1252
rect -4328 1262 -4323 1310
rect -4275 1282 -4270 1290
rect -4247 1282 -4242 1335
rect -4189 1316 -4184 1356
rect -4161 1316 -4156 1356
rect -4141 1334 -4088 1340
rect -4069 1334 -4064 1359
rect -4141 1332 -4096 1334
rect -4088 1327 -4064 1334
rect -4069 1319 -4064 1327
rect -4041 1319 -4036 1359
rect -3960 1343 -3955 1385
rect -3902 1364 -3897 1410
rect -3724 1413 -3720 1418
rect -3649 1413 -3638 1418
rect -3874 1364 -3869 1372
rect -3724 1368 -3719 1413
rect -3643 1395 -3638 1413
rect -3615 1395 -3610 1435
rect -3595 1411 -3590 1419
rect -3328 1418 -3323 1435
rect -3643 1383 -3638 1386
rect -3696 1368 -3691 1376
rect -4021 1335 -3955 1343
rect -4069 1307 -4064 1310
rect -4189 1304 -4184 1307
rect -4328 1245 -4324 1262
rect -4328 1241 -4307 1245
rect -4656 1224 -4651 1227
rect -4628 1224 -4623 1227
rect -4571 1223 -4566 1227
rect -4311 1189 -4307 1241
rect -4275 1234 -4270 1274
rect -4247 1234 -4242 1274
rect -4161 1258 -4156 1307
rect -4227 1250 -4156 1258
rect -4041 1262 -4036 1310
rect -3988 1282 -3983 1290
rect -3960 1282 -3955 1335
rect -3902 1316 -3897 1356
rect -3874 1316 -3869 1356
rect -3854 1332 -3803 1340
rect -3724 1335 -3719 1360
rect -3743 1328 -3719 1335
rect -3724 1320 -3719 1328
rect -3696 1320 -3691 1360
rect -3615 1344 -3610 1386
rect -3557 1365 -3552 1411
rect -3409 1413 -3405 1418
rect -3334 1413 -3323 1418
rect -3529 1365 -3524 1373
rect -3409 1368 -3404 1413
rect -3328 1395 -3323 1413
rect -3300 1395 -3295 1435
rect -3280 1411 -3275 1419
rect -3328 1383 -3323 1386
rect -3381 1368 -3376 1376
rect -3676 1336 -3610 1344
rect -3724 1308 -3719 1311
rect -3902 1304 -3897 1307
rect -4041 1245 -4037 1262
rect -4041 1241 -4020 1245
rect -4275 1222 -4270 1225
rect -4247 1222 -4242 1225
rect -4024 1189 -4020 1241
rect -3988 1234 -3983 1274
rect -3960 1234 -3955 1274
rect -3874 1258 -3869 1307
rect -3940 1250 -3869 1258
rect -3696 1263 -3691 1311
rect -3643 1283 -3638 1291
rect -3615 1283 -3610 1336
rect -3557 1317 -3552 1357
rect -3529 1317 -3524 1357
rect -3509 1335 -3428 1341
rect -3409 1335 -3404 1360
rect -3509 1333 -3436 1335
rect -3428 1328 -3404 1335
rect -3409 1320 -3404 1328
rect -3381 1320 -3376 1360
rect -3300 1344 -3295 1386
rect -3242 1365 -3237 1411
rect -3214 1365 -3209 1373
rect -3361 1336 -3295 1344
rect -3409 1308 -3404 1311
rect -3557 1305 -3552 1308
rect -3696 1246 -3692 1263
rect -3696 1242 -3675 1246
rect -3988 1222 -3983 1225
rect -3960 1222 -3955 1225
rect -3944 1193 -3895 1196
rect -4656 1181 -4651 1189
rect -4628 1181 -4623 1189
rect -4571 1181 -4566 1189
rect -4324 1184 -4307 1189
rect -4037 1184 -4020 1189
rect -4352 1176 -4347 1184
rect -4324 1176 -4319 1184
rect -4267 1176 -4262 1184
rect -4065 1176 -4060 1184
rect -4037 1176 -4032 1184
rect -3980 1176 -3975 1184
rect -4656 1157 -4651 1173
rect -4702 1151 -4651 1157
rect -4656 1133 -4651 1151
rect -4628 1133 -4623 1173
rect -4571 1157 -4566 1173
rect -4608 1149 -4566 1157
rect -4571 1133 -4566 1149
rect -4352 1145 -4347 1168
rect -4375 1138 -4347 1145
rect -4352 1128 -4347 1138
rect -4324 1128 -4319 1168
rect -4267 1152 -4262 1168
rect -4304 1144 -4262 1152
rect -4065 1145 -4060 1168
rect -4267 1128 -4262 1144
rect -4088 1138 -4060 1145
rect -4065 1128 -4060 1138
rect -4037 1128 -4032 1168
rect -3980 1152 -3975 1168
rect -3944 1153 -3940 1193
rect -3899 1183 -3895 1193
rect -3679 1190 -3675 1242
rect -3643 1235 -3638 1275
rect -3615 1235 -3610 1275
rect -3529 1259 -3524 1308
rect -3595 1251 -3524 1259
rect -3381 1263 -3376 1311
rect -3328 1283 -3323 1291
rect -3300 1283 -3295 1336
rect -3242 1317 -3237 1357
rect -3214 1317 -3209 1357
rect -3194 1333 -3186 1341
rect -3242 1305 -3237 1308
rect -3381 1246 -3377 1263
rect -3381 1242 -3360 1246
rect -3643 1223 -3638 1226
rect -3615 1223 -3610 1226
rect -3364 1190 -3360 1242
rect -3328 1235 -3323 1275
rect -3300 1235 -3295 1275
rect -3214 1259 -3209 1308
rect -3280 1251 -3209 1259
rect -3328 1223 -3323 1226
rect -3300 1223 -3295 1226
rect -3285 1194 -3235 1201
rect -3692 1185 -3675 1190
rect -3377 1185 -3360 1190
rect -3899 1180 -3888 1183
rect -3919 1171 -3915 1174
rect -3892 1171 -3888 1180
rect -3720 1177 -3715 1185
rect -3692 1177 -3687 1185
rect -3635 1177 -3630 1185
rect -3405 1177 -3400 1185
rect -3377 1177 -3372 1185
rect -3320 1177 -3315 1185
rect -3844 1171 -3839 1174
rect -4017 1144 -3975 1152
rect -3955 1146 -3940 1153
rect -3919 1144 -3915 1162
rect -3980 1128 -3975 1144
rect -3918 1137 -3915 1144
rect -4656 1121 -4651 1124
rect -4656 1081 -4651 1089
rect -4628 1081 -4623 1124
rect -4571 1120 -4566 1124
rect -3919 1125 -3915 1137
rect -3892 1125 -3888 1162
rect -3844 1142 -3839 1162
rect -3720 1146 -3715 1169
rect -3871 1137 -3839 1142
rect -3743 1139 -3715 1146
rect -3844 1125 -3839 1137
rect -3720 1129 -3715 1139
rect -3692 1129 -3687 1169
rect -3635 1153 -3630 1169
rect -3672 1145 -3630 1153
rect -3405 1146 -3400 1169
rect -3635 1129 -3630 1145
rect -3428 1139 -3400 1146
rect -3405 1129 -3400 1139
rect -3377 1129 -3372 1169
rect -3320 1153 -3315 1169
rect -3285 1154 -3281 1194
rect -3241 1184 -3235 1194
rect -3241 1179 -3228 1184
rect -3259 1172 -3255 1175
rect -3232 1172 -3228 1179
rect -3184 1172 -3179 1175
rect -3357 1145 -3315 1153
rect -3295 1147 -3281 1154
rect -3259 1145 -3255 1163
rect -3320 1129 -3315 1145
rect -3258 1138 -3255 1145
rect -3259 1126 -3255 1138
rect -3232 1126 -3228 1163
rect -3184 1143 -3179 1163
rect -3211 1138 -3179 1143
rect -3184 1126 -3179 1138
rect -4352 1116 -4347 1119
rect -4324 1093 -4319 1119
rect -4267 1115 -4262 1119
rect -4065 1116 -4060 1119
rect -4571 1081 -4566 1089
rect -4037 1092 -4032 1119
rect -3980 1115 -3975 1119
rect -3919 1117 -3915 1120
rect -3892 1116 -3888 1120
rect -3844 1116 -3839 1120
rect -3720 1117 -3715 1120
rect -3692 1090 -3687 1120
rect -3635 1116 -3630 1120
rect -3405 1117 -3400 1120
rect -3377 1097 -3372 1120
rect -3320 1116 -3315 1120
rect -3259 1118 -3255 1121
rect -3232 1117 -3228 1121
rect -3184 1117 -3179 1121
rect -4656 1054 -4651 1073
rect -4693 1048 -4651 1054
rect -4656 1033 -4651 1048
rect -4628 1033 -4623 1073
rect -4571 1057 -4566 1073
rect -4608 1049 -4566 1057
rect -4571 1033 -4566 1049
rect -4275 1026 -4270 1034
rect -4247 1026 -4242 1034
rect -3988 1026 -3983 1034
rect -3960 1026 -3955 1034
rect -3642 1026 -3637 1034
rect -3614 1026 -3609 1034
rect -3360 1026 -3355 1034
rect -3332 1026 -3327 1034
rect -3033 1031 -3028 1039
rect -3005 1031 -3000 1039
rect -4656 1021 -4651 1024
rect -4656 974 -4651 982
rect -4628 974 -4623 1024
rect -4571 1020 -4566 1024
rect -4275 1001 -4270 1018
rect -4356 996 -4352 1001
rect -4281 996 -4270 1001
rect -4571 974 -4566 982
rect -4656 952 -4651 966
rect -4684 946 -4651 952
rect -4656 926 -4651 946
rect -4628 926 -4623 966
rect -4571 950 -4566 966
rect -4356 951 -4351 996
rect -4275 978 -4270 996
rect -4247 978 -4242 1018
rect -4227 994 -4222 1002
rect -3988 1001 -3983 1018
rect -4275 966 -4270 969
rect -4328 951 -4323 959
rect -4608 942 -4566 950
rect -4571 926 -4566 942
rect -4356 918 -4351 943
rect -4656 914 -4651 917
rect -4656 874 -4651 882
rect -4628 874 -4623 917
rect -4571 913 -4566 917
rect -4375 911 -4351 918
rect -4356 903 -4351 911
rect -4328 903 -4323 943
rect -4247 927 -4242 969
rect -4189 948 -4184 994
rect -4069 996 -4065 1001
rect -3994 996 -3983 1001
rect -4161 948 -4156 956
rect -4069 951 -4064 996
rect -3988 978 -3983 996
rect -3960 978 -3955 1018
rect -3940 994 -3935 1002
rect -3642 1001 -3637 1018
rect -3988 966 -3983 969
rect -4041 951 -4036 959
rect -4308 919 -4242 927
rect -4356 891 -4351 894
rect -4571 874 -4566 882
rect -4656 852 -4651 866
rect -4675 846 -4651 852
rect -4656 826 -4651 846
rect -4628 826 -4623 866
rect -4571 850 -4566 866
rect -4608 842 -4566 850
rect -4571 826 -4566 842
rect -4328 846 -4323 894
rect -4275 866 -4270 874
rect -4247 866 -4242 919
rect -4189 900 -4184 940
rect -4161 900 -4156 940
rect -4141 918 -4088 924
rect -4069 918 -4064 943
rect -4141 916 -4096 918
rect -4088 911 -4064 918
rect -4069 903 -4064 911
rect -4041 903 -4036 943
rect -3960 927 -3955 969
rect -3902 948 -3897 994
rect -3723 996 -3719 1001
rect -3648 996 -3637 1001
rect -3874 948 -3869 956
rect -3723 951 -3718 996
rect -3642 978 -3637 996
rect -3614 978 -3609 1018
rect -3594 994 -3589 1002
rect -3360 1001 -3355 1018
rect -3642 966 -3637 969
rect -3695 951 -3690 959
rect -4021 919 -3955 927
rect -4069 891 -4064 894
rect -4189 888 -4184 891
rect -4328 829 -4324 846
rect -4328 825 -4307 829
rect -4656 814 -4651 817
rect -4628 814 -4623 817
rect -4571 813 -4566 817
rect -4311 773 -4307 825
rect -4275 818 -4270 858
rect -4247 818 -4242 858
rect -4161 842 -4156 891
rect -4227 834 -4156 842
rect -4041 846 -4036 894
rect -3988 866 -3983 874
rect -3960 866 -3955 919
rect -3902 900 -3897 940
rect -3874 900 -3869 940
rect -3854 916 -3803 924
rect -3723 918 -3718 943
rect -3742 911 -3718 918
rect -3723 903 -3718 911
rect -3695 903 -3690 943
rect -3614 927 -3609 969
rect -3556 948 -3551 994
rect -3441 996 -3437 1001
rect -3366 996 -3355 1001
rect -3528 948 -3523 956
rect -3441 951 -3436 996
rect -3360 978 -3355 996
rect -3332 978 -3327 1018
rect -3033 1006 -3028 1023
rect -3312 994 -3307 1002
rect -3360 966 -3355 969
rect -3413 951 -3408 959
rect -3675 919 -3609 927
rect -3723 891 -3718 894
rect -3902 888 -3897 891
rect -4041 829 -4037 846
rect -4041 825 -4020 829
rect -4275 806 -4270 809
rect -4247 806 -4242 809
rect -4024 773 -4020 825
rect -3988 818 -3983 858
rect -3960 818 -3955 858
rect -3874 842 -3869 891
rect -3940 834 -3869 842
rect -3695 846 -3690 894
rect -3642 866 -3637 874
rect -3614 866 -3609 919
rect -3556 900 -3551 940
rect -3528 900 -3523 940
rect -3508 918 -3460 924
rect -3441 918 -3436 943
rect -3508 916 -3468 918
rect -3460 911 -3436 918
rect -3441 903 -3436 911
rect -3413 903 -3408 943
rect -3332 927 -3327 969
rect -3274 948 -3269 994
rect -3114 1001 -3110 1006
rect -3039 1001 -3028 1006
rect -3114 956 -3109 1001
rect -3033 983 -3028 1001
rect -3005 983 -3000 1023
rect -2985 999 -2980 1007
rect -3033 971 -3028 974
rect -3086 956 -3081 964
rect -3246 948 -3241 956
rect -3393 919 -3327 927
rect -3441 891 -3436 894
rect -3556 888 -3551 891
rect -3695 829 -3691 846
rect -3695 825 -3674 829
rect -3988 806 -3983 809
rect -3960 806 -3955 809
rect -3945 777 -3895 784
rect -4324 768 -4307 773
rect -4037 768 -4020 773
rect -4657 759 -4652 767
rect -4629 759 -4624 767
rect -4572 759 -4567 767
rect -4352 760 -4347 768
rect -4324 760 -4319 768
rect -4267 760 -4262 768
rect -4065 760 -4060 768
rect -4037 760 -4032 768
rect -3980 760 -3975 768
rect -4657 738 -4652 751
rect -4702 732 -4652 738
rect -4657 711 -4652 732
rect -4629 711 -4624 751
rect -4572 735 -4567 751
rect -4609 727 -4567 735
rect -4352 729 -4347 752
rect -4572 711 -4567 727
rect -4375 722 -4347 729
rect -4352 712 -4347 722
rect -4324 712 -4319 752
rect -4267 736 -4262 752
rect -4304 728 -4262 736
rect -4065 729 -4060 752
rect -4267 712 -4262 728
rect -4088 722 -4060 729
rect -4065 712 -4060 722
rect -4037 712 -4032 752
rect -3980 736 -3975 752
rect -3945 737 -3940 777
rect -3901 767 -3895 777
rect -3678 773 -3674 825
rect -3642 818 -3637 858
rect -3614 818 -3609 858
rect -3528 842 -3523 891
rect -3594 834 -3523 842
rect -3413 846 -3408 894
rect -3360 866 -3355 874
rect -3332 866 -3327 919
rect -3274 900 -3269 940
rect -3246 900 -3241 940
rect -3114 924 -3109 948
rect -3226 916 -3176 924
rect -3133 916 -3109 924
rect -3114 908 -3109 916
rect -3086 908 -3081 948
rect -3005 932 -3000 974
rect -2947 953 -2942 999
rect -2919 953 -2914 961
rect -3066 924 -3000 932
rect -3114 896 -3109 899
rect -3274 888 -3269 891
rect -3413 829 -3409 846
rect -3413 825 -3392 829
rect -3642 806 -3637 809
rect -3614 806 -3609 809
rect -3396 773 -3392 825
rect -3360 818 -3355 858
rect -3332 818 -3327 858
rect -3246 842 -3241 891
rect -3312 834 -3241 842
rect -3086 851 -3081 899
rect -3033 871 -3028 879
rect -3005 871 -3000 924
rect -2947 905 -2942 945
rect -2919 905 -2914 945
rect -2899 921 -2891 929
rect -2947 893 -2942 896
rect -3086 834 -3082 851
rect -3086 830 -3065 834
rect -3360 806 -3355 809
rect -3332 806 -3327 809
rect -3318 778 -3267 785
rect -3069 778 -3065 830
rect -3033 823 -3028 863
rect -3005 823 -3000 863
rect -2919 847 -2914 896
rect -2985 839 -2914 847
rect -3033 811 -3028 814
rect -3005 811 -3000 814
rect -3691 768 -3674 773
rect -3409 768 -3392 773
rect -3901 762 -3888 767
rect -3919 755 -3915 758
rect -3892 755 -3888 762
rect -3719 760 -3714 768
rect -3691 760 -3686 768
rect -3634 760 -3629 768
rect -3437 760 -3432 768
rect -3409 760 -3404 768
rect -3352 760 -3347 768
rect -3844 755 -3839 758
rect -4017 728 -3975 736
rect -3955 730 -3940 737
rect -3919 728 -3915 746
rect -3980 712 -3975 728
rect -3918 721 -3915 728
rect -3919 709 -3915 721
rect -3892 709 -3888 746
rect -3844 726 -3839 746
rect -3719 729 -3714 752
rect -3871 721 -3839 726
rect -3742 722 -3714 729
rect -3844 709 -3839 721
rect -3719 712 -3714 722
rect -3691 712 -3686 752
rect -3634 736 -3629 752
rect -3671 728 -3629 736
rect -3437 729 -3432 752
rect -3634 712 -3629 728
rect -3460 722 -3432 729
rect -3437 712 -3432 722
rect -3409 712 -3404 752
rect -3352 736 -3347 752
rect -3318 737 -3313 778
rect -3273 767 -3267 778
rect -3082 773 -3065 778
rect -3273 762 -3260 767
rect -3110 765 -3105 773
rect -3082 765 -3077 773
rect -3025 765 -3020 773
rect -3291 755 -3287 758
rect -3264 755 -3260 762
rect -3216 755 -3211 758
rect -3389 728 -3347 736
rect -3327 730 -3313 737
rect -3291 728 -3287 746
rect -3352 712 -3347 728
rect -3290 721 -3287 728
rect -4657 699 -4652 702
rect -4657 659 -4652 667
rect -4629 659 -4624 702
rect -4572 698 -4567 702
rect -4352 700 -4347 703
rect -4324 673 -4319 703
rect -4267 699 -4262 703
rect -4065 700 -4060 703
rect -4572 659 -4567 667
rect -4037 671 -4032 703
rect -3980 699 -3975 703
rect -3919 701 -3915 704
rect -3892 700 -3888 704
rect -3844 700 -3839 704
rect -3291 709 -3287 721
rect -3264 709 -3260 746
rect -3216 726 -3211 746
rect -3110 734 -3105 757
rect -3133 727 -3105 734
rect -3243 721 -3211 726
rect -3216 709 -3211 721
rect -3110 717 -3105 727
rect -3082 717 -3077 757
rect -3025 741 -3020 757
rect -3062 733 -3020 741
rect -3025 717 -3020 733
rect -3110 705 -3105 708
rect -3719 700 -3714 703
rect -3691 673 -3686 703
rect -3634 699 -3629 703
rect -3437 700 -3432 703
rect -3409 673 -3404 703
rect -3352 699 -3347 703
rect -3291 701 -3287 704
rect -3264 700 -3260 704
rect -3216 700 -3211 704
rect -3082 686 -3077 708
rect -3025 704 -3020 708
rect -4657 635 -4652 651
rect -4693 629 -4652 635
rect -4657 611 -4652 629
rect -4629 611 -4624 651
rect -4572 635 -4567 651
rect -4609 627 -4567 635
rect -4572 611 -4567 627
rect -4657 599 -4652 602
rect -4657 552 -4652 560
rect -4629 552 -4624 602
rect -4572 598 -4567 602
rect -4275 568 -4270 576
rect -4247 568 -4242 576
rect -3976 568 -3971 576
rect -3948 568 -3943 576
rect -3661 568 -3656 576
rect -3633 568 -3628 576
rect -3332 574 -3327 582
rect -3304 574 -3299 582
rect -3017 574 -3012 582
rect -2989 574 -2984 582
rect -4572 552 -4567 560
rect -4657 533 -4652 544
rect -4684 527 -4652 533
rect -4657 504 -4652 527
rect -4629 504 -4624 544
rect -4572 528 -4567 544
rect -4609 520 -4567 528
rect -4572 504 -4567 520
rect -4657 492 -4652 495
rect -4657 452 -4652 460
rect -4629 452 -4624 495
rect -4572 491 -4567 495
rect -4356 493 -4351 538
rect -4328 493 -4323 548
rect -4275 543 -4270 560
rect -4281 538 -4270 543
rect -4275 520 -4270 538
rect -4247 520 -4242 560
rect -4227 536 -4222 544
rect -3976 543 -3971 560
rect -4275 508 -4270 511
rect -4356 460 -4351 485
rect -4572 452 -4567 460
rect -4375 453 -4351 460
rect -4356 445 -4351 453
rect -4328 445 -4323 485
rect -4247 469 -4242 511
rect -4189 490 -4184 536
rect -3982 538 -3971 543
rect -4161 490 -4156 498
rect -4057 493 -4052 538
rect -3976 520 -3971 538
rect -3948 520 -3943 560
rect -3928 536 -3923 544
rect -3661 543 -3656 560
rect -3976 508 -3971 511
rect -4029 493 -4024 501
rect -4308 461 -4242 469
rect -4657 433 -4652 444
rect -4675 427 -4652 433
rect -4657 404 -4652 427
rect -4629 404 -4624 444
rect -4572 428 -4567 444
rect -4356 433 -4351 436
rect -4609 420 -4567 428
rect -4572 404 -4567 420
rect -4657 392 -4652 395
rect -4629 392 -4624 395
rect -4572 391 -4567 395
rect -4328 388 -4323 436
rect -4275 408 -4270 416
rect -4247 408 -4242 461
rect -4189 442 -4184 482
rect -4161 442 -4156 482
rect -4057 466 -4052 485
rect -4141 458 -4084 466
rect -4076 458 -4052 466
rect -4057 445 -4052 458
rect -4029 445 -4024 485
rect -3948 469 -3943 511
rect -3890 490 -3885 536
rect -3742 538 -3738 543
rect -3667 538 -3656 543
rect -3862 490 -3857 498
rect -3742 493 -3737 538
rect -3661 520 -3656 538
rect -3633 520 -3628 560
rect -3332 549 -3327 566
rect -3413 544 -3409 549
rect -3338 544 -3327 549
rect -3613 536 -3608 544
rect -3661 508 -3656 511
rect -3714 493 -3709 501
rect -4009 461 -3943 469
rect -4057 433 -4052 436
rect -4189 430 -4184 433
rect -4328 371 -4324 388
rect -4328 367 -4307 371
rect -4657 349 -4652 357
rect -4629 349 -4624 357
rect -4572 349 -4567 357
rect -4657 326 -4652 341
rect -4702 320 -4652 326
rect -4657 301 -4652 320
rect -4629 301 -4624 341
rect -4572 325 -4567 341
rect -4609 317 -4567 325
rect -4572 301 -4567 317
rect -4311 315 -4307 367
rect -4275 360 -4270 400
rect -4247 360 -4242 400
rect -4161 384 -4156 433
rect -4227 376 -4156 384
rect -4029 388 -4024 436
rect -3976 408 -3971 416
rect -3948 408 -3943 461
rect -3890 442 -3885 482
rect -3862 442 -3857 482
rect -3842 460 -3761 466
rect -3742 460 -3737 485
rect -3842 458 -3769 460
rect -3761 453 -3737 460
rect -3742 445 -3737 453
rect -3714 445 -3709 485
rect -3633 469 -3628 511
rect -3575 490 -3570 536
rect -3413 499 -3408 544
rect -3332 526 -3327 544
rect -3304 526 -3299 566
rect -3284 542 -3279 550
rect -3017 549 -3012 566
rect -3332 514 -3327 517
rect -3385 499 -3380 507
rect -3547 490 -3542 498
rect -3694 461 -3628 469
rect -3742 433 -3737 436
rect -3890 430 -3885 433
rect -4029 371 -4025 388
rect -4029 367 -4008 371
rect -4275 348 -4270 351
rect -4247 348 -4242 351
rect -4012 315 -4008 367
rect -3976 360 -3971 400
rect -3948 360 -3943 400
rect -3862 384 -3857 433
rect -3928 376 -3857 384
rect -3714 388 -3709 436
rect -3661 408 -3656 416
rect -3633 408 -3628 461
rect -3575 442 -3570 482
rect -3547 442 -3542 482
rect -3413 466 -3408 491
rect -3527 458 -3468 466
rect -3432 459 -3408 466
rect -3413 451 -3408 459
rect -3385 451 -3380 491
rect -3304 475 -3299 517
rect -3246 496 -3241 542
rect -3098 544 -3094 549
rect -3023 544 -3012 549
rect -3218 496 -3213 504
rect -3098 499 -3093 544
rect -3017 526 -3012 544
rect -2989 526 -2984 566
rect -3017 514 -3012 517
rect -3070 499 -3065 507
rect -3365 467 -3299 475
rect -3413 439 -3408 442
rect -3575 430 -3570 433
rect -3714 371 -3710 388
rect -3714 367 -3693 371
rect -3976 348 -3971 351
rect -3948 348 -3943 351
rect -3697 315 -3693 367
rect -3661 360 -3656 400
rect -3633 360 -3628 400
rect -3547 384 -3542 433
rect -3613 376 -3542 384
rect -3385 394 -3380 442
rect -3332 414 -3327 422
rect -3304 414 -3299 467
rect -3246 448 -3241 488
rect -3218 448 -3213 488
rect -3198 466 -3117 472
rect -3098 466 -3093 491
rect -3198 464 -3125 466
rect -3117 459 -3093 466
rect -3098 451 -3093 459
rect -3070 451 -3065 491
rect -2989 475 -2984 517
rect -2931 496 -2926 542
rect -2903 496 -2898 504
rect -3050 467 -2984 475
rect -3098 439 -3093 442
rect -3246 436 -3241 439
rect -3385 377 -3381 394
rect -3385 373 -3364 377
rect -3661 348 -3656 351
rect -3633 348 -3628 351
rect -3368 321 -3364 373
rect -3332 366 -3327 406
rect -3304 366 -3299 406
rect -3218 390 -3213 439
rect -3284 382 -3213 390
rect -3070 394 -3065 442
rect -3017 414 -3012 422
rect -2989 414 -2984 467
rect -2931 448 -2926 488
rect -2903 448 -2898 488
rect -2883 464 -2875 472
rect -2931 436 -2926 439
rect -3070 377 -3066 394
rect -3070 373 -3049 377
rect -3332 354 -3327 357
rect -3304 354 -3299 357
rect -3053 321 -3049 373
rect -3017 366 -3012 406
rect -2989 366 -2984 406
rect -2903 390 -2898 439
rect -2969 382 -2898 390
rect -3017 354 -3012 357
rect -2989 354 -2984 357
rect -3381 316 -3364 321
rect -3066 316 -3049 321
rect -4324 310 -4307 315
rect -4025 310 -4008 315
rect -3710 310 -3693 315
rect -4352 302 -4347 310
rect -4324 302 -4319 310
rect -4267 302 -4262 310
rect -4053 302 -4048 310
rect -4025 302 -4020 310
rect -3968 302 -3963 310
rect -3738 302 -3733 310
rect -3710 302 -3705 310
rect -3653 302 -3648 310
rect -3618 307 -3568 314
rect -3409 308 -3404 316
rect -3381 308 -3376 316
rect -3324 308 -3319 316
rect -3094 308 -3089 316
rect -3066 308 -3061 316
rect -3009 308 -3004 316
rect -2974 313 -2924 320
rect -4657 289 -4652 292
rect -4657 249 -4652 257
rect -4629 249 -4624 292
rect -4572 288 -4567 292
rect -4352 271 -4347 294
rect -4375 264 -4347 271
rect -4572 249 -4567 257
rect -4352 254 -4347 264
rect -4324 254 -4319 294
rect -4267 278 -4262 294
rect -4304 270 -4262 278
rect -4053 271 -4048 294
rect -4267 254 -4262 270
rect -4076 264 -4048 271
rect -4053 254 -4048 264
rect -4025 254 -4020 294
rect -3968 278 -3963 294
rect -4005 270 -3963 278
rect -3738 271 -3733 294
rect -3968 254 -3963 270
rect -3761 264 -3733 271
rect -3738 254 -3733 264
rect -3710 254 -3705 294
rect -3653 278 -3648 294
rect -3618 279 -3613 307
rect -3574 289 -3568 307
rect -3574 284 -3561 289
rect -3690 270 -3648 278
rect -3628 272 -3613 279
rect -3592 277 -3588 280
rect -3565 277 -3561 284
rect -3517 277 -3512 280
rect -3409 277 -3404 300
rect -3653 254 -3648 270
rect -3432 270 -3404 277
rect -3592 250 -3588 268
rect -4352 242 -4347 245
rect -4324 242 -4319 245
rect -4267 241 -4262 245
rect -4053 242 -4048 245
rect -4657 223 -4652 241
rect -4693 217 -4652 223
rect -4657 201 -4652 217
rect -4629 201 -4624 241
rect -4572 225 -4567 241
rect -4609 217 -4567 225
rect -4025 225 -4020 245
rect -3968 241 -3963 245
rect -3738 242 -3733 245
rect -4572 201 -4567 217
rect -3710 207 -3705 245
rect -3653 241 -3648 245
rect -3591 243 -3588 250
rect -3592 231 -3588 243
rect -3565 231 -3561 268
rect -3517 248 -3512 268
rect -3409 260 -3404 270
rect -3381 260 -3376 300
rect -3324 284 -3319 300
rect -3361 276 -3319 284
rect -3094 277 -3089 300
rect -3324 260 -3319 276
rect -3117 270 -3089 277
rect -3094 260 -3089 270
rect -3066 260 -3061 300
rect -3009 284 -3004 300
rect -2974 285 -2969 313
rect -2930 295 -2924 313
rect -2930 290 -2917 295
rect -3046 276 -3004 284
rect -2984 278 -2969 285
rect -2948 283 -2944 286
rect -2921 283 -2917 290
rect -2873 283 -2868 286
rect -3009 260 -3004 276
rect -2948 256 -2944 274
rect -3409 248 -3404 251
rect -3544 243 -3512 248
rect -3517 231 -3512 243
rect -3592 223 -3588 226
rect -3565 222 -3561 226
rect -3517 222 -3512 226
rect -3381 221 -3376 251
rect -3324 247 -3319 251
rect -3094 248 -3089 251
rect -3066 211 -3061 251
rect -3009 247 -3004 251
rect -2947 249 -2944 256
rect -2948 237 -2944 249
rect -2921 237 -2917 274
rect -2873 254 -2868 274
rect -2900 249 -2868 254
rect -2873 237 -2868 249
rect -2948 229 -2944 232
rect -2921 228 -2917 232
rect -2873 228 -2868 232
rect -4275 194 -4270 202
rect -4247 194 -4242 202
rect -4657 189 -4652 192
rect -4657 142 -4652 150
rect -4629 142 -4624 192
rect -4572 188 -4567 192
rect -4356 164 -4352 169
rect -4572 142 -4567 150
rect -4657 121 -4652 134
rect -4684 115 -4652 121
rect -4657 94 -4652 115
rect -4629 94 -4624 134
rect -4572 118 -4567 134
rect -4356 119 -4351 164
rect -4328 119 -4323 172
rect -4275 169 -4270 186
rect -4281 164 -4270 169
rect -4275 146 -4270 164
rect -4247 146 -4242 186
rect -4227 162 -4222 170
rect -4275 134 -4270 137
rect -4609 110 -4567 118
rect -4572 94 -4567 110
rect -4356 86 -4351 111
rect -4657 82 -4652 85
rect -4657 42 -4652 50
rect -4629 42 -4624 85
rect -4572 81 -4567 85
rect -4375 79 -4351 86
rect -4356 71 -4351 79
rect -4328 71 -4323 111
rect -4247 95 -4242 137
rect -4189 116 -4184 162
rect -3944 161 -3939 169
rect -3916 161 -3911 169
rect -3629 161 -3624 169
rect -3601 161 -3596 169
rect -3944 136 -3939 153
rect -4025 131 -4021 136
rect -3950 131 -3939 136
rect -4161 116 -4156 124
rect -4308 87 -4242 95
rect -4356 59 -4351 62
rect -4572 42 -4567 50
rect -4657 21 -4652 34
rect -4675 15 -4652 21
rect -4657 -6 -4652 15
rect -4629 -6 -4624 34
rect -4572 18 -4567 34
rect -4609 10 -4567 18
rect -4572 -6 -4567 10
rect -4328 14 -4323 62
rect -4275 34 -4270 42
rect -4247 34 -4242 87
rect -4189 68 -4184 108
rect -4161 68 -4156 108
rect -4025 86 -4020 131
rect -3944 113 -3939 131
rect -3916 113 -3911 153
rect -3896 129 -3891 137
rect -3629 136 -3624 153
rect -3944 101 -3939 104
rect -3997 86 -3992 94
rect -4189 56 -4184 59
rect -4328 -3 -4324 14
rect -4328 -7 -4307 -3
rect -4657 -18 -4652 -15
rect -4629 -18 -4624 -15
rect -4572 -19 -4567 -15
rect -4311 -59 -4307 -7
rect -4275 -14 -4270 26
rect -4247 -14 -4242 26
rect -4161 10 -4156 59
rect -4025 53 -4020 78
rect -4044 46 -4020 53
rect -4025 38 -4020 46
rect -3997 38 -3992 78
rect -3916 62 -3911 104
rect -3858 83 -3853 129
rect -3710 131 -3706 136
rect -3635 131 -3624 136
rect -3830 83 -3825 91
rect -3710 86 -3705 131
rect -3629 113 -3624 131
rect -3601 113 -3596 153
rect -3581 129 -3576 137
rect -3629 101 -3624 104
rect -3682 86 -3677 94
rect -3977 54 -3911 62
rect -4025 26 -4020 29
rect -4227 2 -4156 10
rect -3997 -19 -3992 29
rect -3944 1 -3939 9
rect -3916 1 -3911 54
rect -3858 35 -3853 75
rect -3830 35 -3825 75
rect -3810 53 -3729 59
rect -3710 53 -3705 78
rect -3810 51 -3737 53
rect -3729 46 -3705 53
rect -3710 38 -3705 46
rect -3682 38 -3677 78
rect -3601 62 -3596 104
rect -3543 83 -3538 129
rect -3515 83 -3510 91
rect -3662 54 -3596 62
rect -3710 26 -3705 29
rect -3858 23 -3853 26
rect -4275 -26 -4270 -23
rect -4247 -26 -4242 -23
rect -3997 -36 -3993 -19
rect -3997 -40 -3976 -36
rect -4324 -64 -4307 -59
rect -4352 -72 -4347 -64
rect -4324 -72 -4319 -64
rect -4267 -72 -4262 -64
rect -4352 -103 -4347 -80
rect -4375 -110 -4347 -103
rect -4352 -120 -4347 -110
rect -4324 -120 -4319 -80
rect -4267 -96 -4262 -80
rect -3980 -92 -3976 -40
rect -3944 -47 -3939 -7
rect -3916 -47 -3911 -7
rect -3830 -23 -3825 26
rect -3896 -31 -3825 -23
rect -3682 -19 -3677 29
rect -3629 1 -3624 9
rect -3601 1 -3596 54
rect -3543 35 -3538 75
rect -3515 35 -3510 75
rect -3495 51 -3487 59
rect -3543 23 -3538 26
rect -3682 -36 -3678 -19
rect -3682 -40 -3661 -36
rect -3944 -59 -3939 -56
rect -3916 -59 -3911 -56
rect -3665 -92 -3661 -40
rect -3629 -47 -3624 -7
rect -3601 -47 -3596 -7
rect -3515 -23 -3510 26
rect -3581 -31 -3510 -23
rect -3629 -59 -3624 -56
rect -3601 -59 -3596 -56
rect -4304 -104 -4262 -96
rect -3993 -97 -3976 -92
rect -3678 -97 -3661 -92
rect -4267 -120 -4262 -104
rect -4021 -105 -4016 -97
rect -3993 -105 -3988 -97
rect -3936 -105 -3931 -97
rect -3706 -105 -3701 -97
rect -3678 -105 -3673 -97
rect -3621 -105 -3616 -97
rect -3586 -100 -3536 -93
rect -4352 -132 -4347 -129
rect -4324 -132 -4319 -129
rect -4267 -133 -4262 -129
rect -4021 -136 -4016 -113
rect -4044 -143 -4016 -136
rect -4021 -153 -4016 -143
rect -3993 -153 -3988 -113
rect -3936 -129 -3931 -113
rect -3973 -137 -3931 -129
rect -3706 -136 -3701 -113
rect -3936 -153 -3931 -137
rect -3729 -143 -3701 -136
rect -3706 -153 -3701 -143
rect -3678 -153 -3673 -113
rect -3621 -129 -3616 -113
rect -3586 -128 -3581 -100
rect -3542 -118 -3536 -100
rect -3542 -123 -3529 -118
rect -3658 -137 -3616 -129
rect -3596 -135 -3581 -128
rect -3560 -130 -3556 -127
rect -3533 -130 -3529 -123
rect -3485 -130 -3480 -127
rect -3621 -153 -3616 -137
rect -3560 -157 -3556 -139
rect -4021 -165 -4016 -162
rect -4275 -182 -4270 -174
rect -4247 -182 -4242 -174
rect -4356 -212 -4352 -207
rect -4356 -257 -4351 -212
rect -4328 -257 -4323 -199
rect -4275 -207 -4270 -190
rect -4281 -212 -4270 -207
rect -4275 -230 -4270 -212
rect -4247 -230 -4242 -190
rect -3993 -192 -3988 -162
rect -3936 -166 -3931 -162
rect -3706 -165 -3701 -162
rect -3678 -201 -3673 -162
rect -3621 -166 -3616 -162
rect -3559 -164 -3556 -157
rect -3560 -176 -3556 -164
rect -3533 -176 -3529 -139
rect -3485 -159 -3480 -139
rect -3512 -164 -3480 -159
rect -3485 -176 -3480 -164
rect -3560 -184 -3556 -181
rect -3533 -185 -3529 -181
rect -3485 -185 -3480 -181
rect -4227 -214 -4222 -206
rect -4275 -242 -4270 -239
rect -4356 -290 -4351 -265
rect -4375 -297 -4351 -290
rect -4356 -305 -4351 -297
rect -4328 -305 -4323 -265
rect -4247 -281 -4242 -239
rect -4189 -260 -4184 -214
rect -4161 -260 -4156 -252
rect -4308 -289 -4242 -281
rect -4356 -317 -4351 -314
rect -4328 -362 -4323 -314
rect -4275 -342 -4270 -334
rect -4247 -342 -4242 -289
rect -4189 -308 -4184 -268
rect -4161 -308 -4156 -268
rect -4141 -292 -4133 -284
rect -4189 -320 -4184 -317
rect -4328 -379 -4324 -362
rect -4328 -383 -4307 -379
rect -4311 -435 -4307 -383
rect -4275 -390 -4270 -350
rect -4247 -390 -4242 -350
rect -4161 -366 -4156 -317
rect -4227 -374 -4156 -366
rect -4275 -402 -4270 -399
rect -4247 -402 -4242 -399
rect -4324 -440 -4307 -435
rect -4352 -448 -4347 -440
rect -4324 -448 -4319 -440
rect -4267 -448 -4262 -440
rect -4352 -479 -4347 -456
rect -4375 -486 -4347 -479
rect -4352 -496 -4347 -486
rect -4324 -496 -4319 -456
rect -4267 -472 -4262 -456
rect -4304 -480 -4262 -472
rect -4267 -496 -4262 -480
rect -4352 -508 -4347 -505
rect -4324 -508 -4319 -505
rect -4267 -509 -4262 -505
<< polycontact >>
rect -4708 1553 -4702 1559
rect -4616 1559 -4608 1567
rect -4699 1450 -4693 1456
rect -4616 1459 -4608 1467
rect -4352 1412 -4348 1417
rect -4285 1412 -4281 1417
rect -4690 1348 -4684 1354
rect -4235 1410 -4227 1418
rect -4222 1410 -4215 1418
rect -4190 1410 -4184 1418
rect -4616 1352 -4608 1360
rect -4383 1327 -4375 1334
rect -4065 1412 -4061 1417
rect -3998 1412 -3994 1417
rect -3948 1410 -3940 1418
rect -3935 1410 -3928 1418
rect -3903 1410 -3897 1418
rect -4316 1335 -4308 1343
rect -4681 1248 -4675 1254
rect -4616 1252 -4608 1260
rect -4149 1332 -4141 1340
rect -4096 1327 -4088 1334
rect -3720 1413 -3716 1418
rect -3653 1413 -3649 1418
rect -3603 1411 -3595 1419
rect -3590 1411 -3583 1419
rect -3558 1411 -3552 1419
rect -4029 1335 -4021 1343
rect -4324 1256 -4319 1262
rect -4280 1256 -4275 1262
rect -4235 1250 -4227 1258
rect -3862 1332 -3854 1340
rect -3803 1332 -3795 1340
rect -3751 1328 -3743 1335
rect -3405 1413 -3401 1418
rect -3338 1413 -3334 1418
rect -3288 1411 -3280 1419
rect -3275 1411 -3268 1419
rect -3243 1411 -3237 1419
rect -3684 1336 -3676 1344
rect -4037 1256 -4032 1262
rect -3993 1256 -3988 1262
rect -3948 1250 -3940 1258
rect -3517 1333 -3509 1341
rect -3436 1328 -3428 1335
rect -3369 1336 -3361 1344
rect -3692 1257 -3687 1263
rect -3648 1257 -3643 1263
rect -4708 1151 -4702 1157
rect -4616 1149 -4608 1157
rect -4383 1138 -4375 1145
rect -4312 1144 -4304 1152
rect -4096 1138 -4088 1145
rect -3603 1251 -3595 1259
rect -3202 1333 -3194 1341
rect -3377 1257 -3372 1263
rect -3333 1257 -3328 1263
rect -3288 1251 -3280 1259
rect -4025 1144 -4017 1152
rect -3960 1146 -3955 1153
rect -3925 1137 -3918 1144
rect -3876 1137 -3871 1142
rect -3751 1139 -3743 1146
rect -3680 1145 -3672 1153
rect -3436 1139 -3428 1146
rect -3365 1145 -3357 1153
rect -3300 1147 -3295 1154
rect -3265 1138 -3258 1145
rect -3216 1138 -3211 1143
rect -4324 1086 -4319 1093
rect -4037 1088 -4032 1092
rect -3377 1092 -3372 1097
rect -3692 1086 -3687 1090
rect -4699 1048 -4693 1054
rect -4616 1049 -4608 1057
rect -4352 996 -4348 1001
rect -4285 996 -4281 1001
rect -4690 946 -4684 952
rect -4235 994 -4227 1002
rect -4222 994 -4215 1002
rect -4190 994 -4184 1002
rect -4616 942 -4608 950
rect -4383 911 -4375 918
rect -4065 996 -4061 1001
rect -3998 996 -3994 1001
rect -3948 994 -3940 1002
rect -3935 994 -3928 1002
rect -3903 994 -3897 1002
rect -4316 919 -4308 927
rect -4681 846 -4675 852
rect -4616 842 -4608 850
rect -4149 916 -4141 924
rect -4096 911 -4088 918
rect -3719 996 -3715 1001
rect -3652 996 -3648 1001
rect -3602 994 -3594 1002
rect -3589 994 -3582 1002
rect -3557 994 -3551 1002
rect -4029 919 -4021 927
rect -4324 840 -4319 846
rect -4280 840 -4275 846
rect -4235 834 -4227 842
rect -3862 916 -3854 924
rect -3803 916 -3796 924
rect -3750 911 -3742 918
rect -3437 996 -3433 1001
rect -3370 996 -3366 1001
rect -3320 994 -3312 1002
rect -3307 994 -3300 1002
rect -3275 994 -3269 1002
rect -3683 919 -3675 927
rect -4037 840 -4032 846
rect -3993 840 -3988 846
rect -3948 834 -3940 842
rect -3516 916 -3508 924
rect -3468 911 -3460 918
rect -3110 1001 -3106 1006
rect -3043 1001 -3039 1006
rect -2993 999 -2985 1007
rect -2980 999 -2973 1007
rect -2948 999 -2942 1007
rect -3401 919 -3393 927
rect -3691 840 -3686 846
rect -3647 840 -3642 846
rect -4708 732 -4702 738
rect -4617 727 -4609 735
rect -4383 722 -4375 729
rect -4312 728 -4304 736
rect -4096 722 -4088 729
rect -3602 834 -3594 842
rect -3234 916 -3226 924
rect -3176 916 -3169 924
rect -3141 916 -3133 924
rect -3074 924 -3066 932
rect -3409 840 -3404 846
rect -3365 840 -3360 846
rect -3320 834 -3312 842
rect -2907 921 -2899 929
rect -3082 845 -3077 851
rect -3038 845 -3033 851
rect -2993 839 -2985 847
rect -4025 728 -4017 736
rect -3960 730 -3955 737
rect -3925 721 -3918 728
rect -3876 721 -3871 726
rect -3750 722 -3742 729
rect -3679 728 -3671 736
rect -3468 722 -3460 729
rect -3397 728 -3389 736
rect -3332 730 -3327 737
rect -3297 721 -3290 728
rect -4324 666 -4319 673
rect -3141 727 -3133 734
rect -3248 721 -3243 726
rect -3070 733 -3062 741
rect -4037 663 -4032 671
rect -3691 669 -3686 673
rect -3082 679 -3077 686
rect -3409 665 -3404 673
rect -4699 629 -4693 635
rect -4617 627 -4609 635
rect -4328 548 -4323 555
rect -4690 527 -4684 533
rect -4617 520 -4609 528
rect -4356 538 -4351 543
rect -4285 538 -4281 543
rect -4235 536 -4227 544
rect -4222 536 -4215 544
rect -4190 536 -4184 544
rect -4383 453 -4375 460
rect -4057 538 -4052 543
rect -3986 538 -3982 543
rect -3936 536 -3928 544
rect -3923 536 -3916 544
rect -3891 536 -3885 544
rect -4316 461 -4308 469
rect -4681 427 -4675 433
rect -4617 420 -4609 428
rect -4149 458 -4141 466
rect -4084 458 -4076 466
rect -3738 538 -3734 543
rect -3671 538 -3667 543
rect -3409 544 -3405 549
rect -3342 544 -3338 549
rect -3621 536 -3613 544
rect -3608 536 -3601 544
rect -3576 536 -3570 544
rect -4017 461 -4009 469
rect -4324 382 -4319 388
rect -4280 382 -4275 388
rect -4708 320 -4702 326
rect -4617 317 -4609 325
rect -4235 376 -4227 384
rect -3850 458 -3842 466
rect -3769 453 -3761 460
rect -3292 542 -3284 550
rect -3279 542 -3272 550
rect -3247 542 -3241 550
rect -3702 461 -3694 469
rect -4025 382 -4020 388
rect -3981 382 -3976 388
rect -3936 376 -3928 384
rect -3535 458 -3527 466
rect -3468 458 -3460 466
rect -3440 459 -3432 466
rect -3094 544 -3090 549
rect -3027 544 -3023 549
rect -2932 542 -2926 550
rect -3373 467 -3365 475
rect -3710 382 -3705 388
rect -3666 382 -3661 388
rect -3621 376 -3613 384
rect -3206 464 -3198 472
rect -3125 459 -3117 466
rect -3058 467 -3050 475
rect -3381 388 -3376 394
rect -3337 388 -3332 394
rect -3292 382 -3284 390
rect -2891 464 -2883 472
rect -3066 388 -3061 394
rect -3022 388 -3017 394
rect -2977 382 -2969 390
rect -4383 264 -4375 271
rect -4312 270 -4304 278
rect -4084 264 -4076 271
rect -4013 270 -4005 278
rect -3769 264 -3761 271
rect -3698 270 -3690 278
rect -3633 272 -3628 279
rect -3440 270 -3432 277
rect -4699 217 -4693 223
rect -4617 217 -4609 225
rect -4025 219 -4020 225
rect -3598 243 -3591 250
rect -3369 276 -3361 284
rect -3125 270 -3117 277
rect -3054 276 -3046 284
rect -2989 278 -2984 285
rect -3549 243 -3544 248
rect -3381 217 -3376 221
rect -2954 249 -2947 256
rect -2905 249 -2900 254
rect -3710 199 -3705 207
rect -3066 206 -3061 211
rect -4328 172 -4323 178
rect -4352 164 -4348 169
rect -4690 115 -4684 121
rect -4285 164 -4281 169
rect -4235 162 -4227 170
rect -4222 162 -4215 170
rect -4190 162 -4184 170
rect -4617 110 -4609 118
rect -4383 79 -4375 86
rect -4021 131 -4017 136
rect -3954 131 -3950 136
rect -4316 87 -4308 95
rect -4681 15 -4675 21
rect -4617 10 -4609 18
rect -4149 84 -4141 92
rect -3904 129 -3896 137
rect -3891 129 -3884 137
rect -3859 129 -3853 137
rect -4324 8 -4319 14
rect -4280 8 -4275 14
rect -4052 46 -4044 53
rect -3706 131 -3702 136
rect -3639 131 -3635 136
rect -3589 129 -3581 137
rect -3576 129 -3569 137
rect -3544 129 -3538 137
rect -3985 54 -3977 62
rect -4235 2 -4227 10
rect -3818 51 -3810 59
rect -3737 46 -3729 53
rect -3670 54 -3662 62
rect -3993 -25 -3988 -19
rect -3949 -25 -3944 -19
rect -4383 -110 -4375 -103
rect -3904 -31 -3896 -23
rect -3503 51 -3495 59
rect -3678 -25 -3673 -19
rect -3634 -25 -3629 -19
rect -3589 -31 -3581 -23
rect -4312 -104 -4304 -96
rect -4052 -143 -4044 -136
rect -3981 -137 -3973 -129
rect -3737 -143 -3729 -136
rect -3666 -137 -3658 -129
rect -3601 -135 -3596 -128
rect -4328 -199 -4323 -194
rect -4352 -212 -4348 -207
rect -4285 -212 -4281 -207
rect -3993 -199 -3988 -192
rect -3566 -164 -3559 -157
rect -3517 -164 -3512 -159
rect -3678 -205 -3673 -201
rect -4235 -214 -4227 -206
rect -4222 -214 -4215 -206
rect -4190 -214 -4184 -206
rect -4383 -297 -4375 -290
rect -4316 -289 -4308 -281
rect -4149 -292 -4141 -284
rect -4324 -368 -4319 -362
rect -4280 -368 -4275 -362
rect -4235 -374 -4227 -366
rect -4383 -486 -4375 -479
rect -4312 -480 -4304 -472
<< metal1 >>
rect -4665 1606 -4646 1612
rect -4639 1606 -4622 1612
rect -4615 1606 -4573 1612
rect -4565 1606 -4555 1612
rect -4546 1606 -4541 1612
rect -4665 1591 -4658 1606
rect -4616 1591 -4609 1606
rect -4580 1591 -4573 1606
rect -4643 1567 -4636 1583
rect -4558 1572 -4551 1583
rect -4643 1559 -4616 1567
rect -4708 1157 -4702 1553
rect -4616 1543 -4608 1559
rect -4558 1558 -4552 1572
rect -4558 1554 -4551 1558
rect -4424 1554 -4418 1621
rect -4558 1548 -4418 1554
rect -4558 1543 -4551 1548
rect -4670 1525 -4662 1534
rect -4587 1525 -4579 1534
rect -4662 1517 -4658 1525
rect -4650 1517 -4622 1525
rect -4614 1517 -4579 1525
rect -4570 1517 -4560 1525
rect -4551 1522 -4550 1525
rect -4425 1524 -4417 1528
rect -4551 1517 -4446 1522
rect -4665 1506 -4646 1512
rect -4639 1506 -4619 1512
rect -4611 1506 -4573 1512
rect -4565 1506 -4555 1512
rect -4546 1506 -4541 1512
rect -4665 1491 -4658 1506
rect -4616 1491 -4609 1506
rect -4580 1491 -4573 1506
rect -4454 1503 -4446 1517
rect -4454 1495 -4376 1503
rect -4643 1467 -4636 1483
rect -4643 1459 -4616 1467
rect -4708 738 -4702 1151
rect -4708 326 -4702 732
rect -4699 1054 -4693 1450
rect -4616 1443 -4608 1459
rect -4558 1465 -4551 1483
rect -4558 1457 -4496 1465
rect -4278 1457 -4265 1464
rect -4258 1457 -4244 1464
rect -4237 1457 -4225 1464
rect -3991 1457 -3978 1464
rect -3971 1457 -3957 1464
rect -3950 1457 -3938 1464
rect -3646 1458 -3633 1465
rect -3626 1458 -3612 1465
rect -3605 1458 -3593 1465
rect -3331 1458 -3318 1465
rect -3311 1458 -3297 1465
rect -3290 1458 -3278 1465
rect -4558 1443 -4551 1457
rect -4284 1442 -4277 1457
rect -4235 1442 -4228 1457
rect -3997 1442 -3990 1457
rect -3948 1442 -3941 1457
rect -3652 1443 -3645 1458
rect -3603 1443 -3596 1458
rect -3337 1443 -3330 1458
rect -3288 1443 -3281 1458
rect -4670 1425 -4662 1434
rect -4587 1425 -4579 1434
rect -4662 1417 -4658 1425
rect -4650 1417 -4622 1425
rect -4614 1417 -4579 1425
rect -4570 1417 -4560 1425
rect -4551 1417 -4550 1425
rect -4262 1418 -4255 1434
rect -3975 1418 -3968 1434
rect -3630 1419 -3623 1435
rect -3315 1419 -3308 1435
rect -4348 1412 -4285 1417
rect -4262 1410 -4235 1418
rect -4215 1410 -4190 1418
rect -4061 1412 -3998 1417
rect -3975 1410 -3948 1418
rect -3928 1410 -3903 1418
rect -3716 1413 -3653 1418
rect -3630 1411 -3603 1419
rect -3583 1411 -3558 1419
rect -3401 1413 -3338 1418
rect -3315 1411 -3288 1419
rect -3268 1411 -3243 1419
rect -4665 1399 -4646 1405
rect -4639 1399 -4573 1405
rect -4565 1399 -4555 1405
rect -4546 1399 -4541 1405
rect -4536 1399 -4360 1405
rect -4665 1384 -4658 1399
rect -4616 1384 -4609 1399
rect -4580 1384 -4573 1399
rect -4537 1398 -4360 1399
rect -4366 1389 -4360 1398
rect -4235 1394 -4227 1410
rect -3948 1394 -3940 1410
rect -3603 1395 -3595 1411
rect -3288 1395 -3280 1411
rect -4366 1382 -4365 1389
rect -4360 1382 -4346 1389
rect -4339 1382 -4325 1389
rect -4318 1382 -4304 1389
rect -4643 1360 -4636 1376
rect -4699 635 -4693 1048
rect -4699 223 -4693 629
rect -4643 1352 -4616 1360
rect -4690 952 -4684 1348
rect -4616 1336 -4608 1352
rect -4558 1358 -4551 1376
rect -4365 1367 -4358 1382
rect -4316 1367 -4309 1382
rect -4289 1376 -4281 1385
rect -4191 1381 -4179 1386
rect -4198 1379 -4179 1381
rect -4172 1379 -4158 1386
rect -4151 1379 -4133 1386
rect -4073 1382 -4059 1389
rect -4052 1382 -4038 1389
rect -4031 1382 -4017 1389
rect -4289 1368 -4277 1376
rect -4269 1368 -4224 1376
rect -4198 1364 -4191 1379
rect -4149 1364 -4142 1379
rect -4558 1350 -4508 1358
rect -4558 1336 -4551 1350
rect -4343 1343 -4336 1359
rect -4078 1367 -4071 1382
rect -4029 1367 -4022 1382
rect -4002 1376 -3994 1385
rect -3904 1381 -3892 1386
rect -3911 1379 -3892 1381
rect -3885 1379 -3871 1386
rect -3864 1383 -3733 1386
rect -3728 1383 -3714 1390
rect -3707 1383 -3693 1390
rect -3686 1383 -3672 1390
rect -3864 1379 -3726 1383
rect -4002 1368 -3990 1376
rect -3982 1368 -3937 1376
rect -3911 1364 -3904 1379
rect -3862 1364 -3855 1379
rect -4343 1335 -4316 1343
rect -4670 1318 -4662 1327
rect -4587 1318 -4579 1327
rect -4662 1310 -4658 1318
rect -4650 1310 -4622 1318
rect -4614 1310 -4579 1318
rect -4570 1310 -4560 1318
rect -4551 1310 -4550 1318
rect -4665 1299 -4646 1305
rect -4639 1299 -4619 1305
rect -4612 1299 -4573 1305
rect -4565 1299 -4555 1305
rect -4546 1299 -4541 1305
rect -4665 1284 -4658 1299
rect -4616 1284 -4609 1299
rect -4580 1284 -4573 1299
rect -4643 1260 -4636 1276
rect -4690 533 -4684 946
rect -4690 121 -4684 527
rect -4643 1252 -4616 1260
rect -4681 852 -4675 1248
rect -4616 1236 -4608 1252
rect -4558 1257 -4551 1276
rect -4558 1250 -4530 1257
rect -4558 1236 -4551 1250
rect -4670 1218 -4662 1227
rect -4587 1218 -4579 1227
rect -4662 1210 -4658 1218
rect -4650 1210 -4622 1218
rect -4614 1210 -4579 1218
rect -4570 1210 -4560 1218
rect -4551 1210 -4550 1218
rect -4665 1196 -4646 1202
rect -4639 1196 -4623 1202
rect -4616 1196 -4573 1202
rect -4565 1196 -4555 1202
rect -4546 1196 -4541 1202
rect -4665 1181 -4658 1196
rect -4616 1181 -4609 1196
rect -4580 1181 -4573 1196
rect -4643 1157 -4636 1173
rect -4643 1149 -4616 1157
rect -4616 1133 -4608 1149
rect -4558 1154 -4551 1173
rect -4383 1154 -4375 1327
rect -4316 1319 -4308 1335
rect -4176 1340 -4169 1356
rect -4056 1343 -4049 1359
rect -4176 1332 -4149 1340
rect -4056 1335 -4029 1343
rect -4149 1316 -4141 1332
rect -4370 1301 -4362 1310
rect -4364 1293 -4358 1301
rect -4350 1293 -4300 1301
rect -4278 1297 -4265 1304
rect -4258 1297 -4241 1304
rect -4234 1297 -4219 1304
rect -4203 1298 -4195 1307
rect -4284 1282 -4277 1297
rect -4235 1282 -4228 1297
rect -4194 1290 -4191 1298
rect -4183 1290 -4133 1298
rect -4319 1256 -4280 1262
rect -4262 1258 -4255 1274
rect -4262 1250 -4235 1258
rect -4235 1234 -4227 1250
rect -4289 1217 -4281 1225
rect -4281 1208 -4277 1216
rect -4269 1208 -4249 1216
rect -4241 1208 -4225 1216
rect -4356 1191 -4342 1197
rect -4335 1191 -4321 1197
rect -4314 1191 -4269 1197
rect -4261 1191 -4251 1197
rect -4242 1191 -4239 1197
rect -4356 1190 -4354 1191
rect -4361 1176 -4354 1190
rect -4312 1176 -4305 1191
rect -4276 1176 -4269 1191
rect -4558 1147 -4375 1154
rect -4558 1133 -4551 1147
rect -4383 1145 -4375 1147
rect -4339 1152 -4332 1168
rect -4254 1153 -4247 1168
rect -4339 1144 -4312 1152
rect -4312 1128 -4304 1144
rect -4254 1128 -4247 1145
rect -4670 1115 -4662 1124
rect -4587 1115 -4579 1124
rect -4366 1115 -4358 1119
rect -4662 1107 -4658 1115
rect -4650 1107 -4622 1115
rect -4614 1107 -4579 1115
rect -4570 1107 -4560 1115
rect -4551 1110 -4358 1115
rect -4283 1110 -4275 1119
rect -4236 1111 -4227 1208
rect -4096 1145 -4088 1327
rect -4029 1319 -4021 1335
rect -3889 1340 -3882 1356
rect -3889 1332 -3862 1340
rect -3862 1316 -3854 1332
rect -4083 1301 -4075 1310
rect -4077 1293 -4071 1301
rect -4063 1293 -4013 1301
rect -3991 1297 -3978 1304
rect -3971 1297 -3954 1304
rect -3947 1297 -3932 1304
rect -3916 1298 -3908 1307
rect -3997 1282 -3990 1297
rect -3948 1282 -3941 1297
rect -3907 1290 -3904 1298
rect -3896 1290 -3846 1298
rect -4032 1256 -3993 1262
rect -3975 1258 -3968 1274
rect -3975 1250 -3948 1258
rect -3948 1234 -3940 1250
rect -4002 1217 -3994 1225
rect -3994 1208 -3990 1216
rect -3982 1208 -3962 1216
rect -3954 1208 -3938 1216
rect -4069 1191 -4055 1197
rect -4048 1191 -4034 1197
rect -4027 1191 -3982 1197
rect -3974 1191 -3964 1197
rect -3955 1191 -3952 1197
rect -4069 1190 -4067 1191
rect -4074 1176 -4067 1190
rect -4025 1176 -4018 1191
rect -3989 1176 -3982 1191
rect -4052 1152 -4045 1168
rect -4052 1144 -4025 1152
rect -4025 1128 -4017 1144
rect -3967 1128 -3960 1168
rect -4079 1111 -4071 1119
rect -4236 1110 -4071 1111
rect -3996 1110 -3988 1119
rect -3949 1110 -3940 1208
rect -3839 1192 -3834 1379
rect -3733 1368 -3726 1379
rect -3684 1368 -3677 1383
rect -3657 1377 -3649 1386
rect -3559 1382 -3547 1387
rect -3566 1380 -3547 1382
rect -3540 1380 -3526 1387
rect -3519 1380 -3501 1387
rect -3413 1383 -3399 1390
rect -3392 1383 -3378 1390
rect -3371 1383 -3357 1390
rect -3657 1369 -3645 1377
rect -3637 1369 -3592 1377
rect -3566 1365 -3559 1380
rect -3517 1365 -3510 1380
rect -3711 1344 -3704 1360
rect -3418 1368 -3411 1383
rect -3369 1368 -3362 1383
rect -3342 1377 -3334 1386
rect -3244 1382 -3232 1387
rect -3251 1380 -3232 1382
rect -3225 1380 -3211 1387
rect -3204 1380 -3174 1387
rect -3342 1369 -3330 1377
rect -3322 1369 -3277 1377
rect -3251 1365 -3244 1380
rect -3202 1365 -3195 1380
rect -3795 1332 -3781 1340
rect -3711 1336 -3684 1344
rect -3927 1186 -3918 1192
rect -3912 1186 -3892 1192
rect -3886 1186 -3865 1192
rect -3859 1186 -3846 1192
rect -3840 1186 -3834 1192
rect -3927 1171 -3922 1186
rect -3854 1171 -3849 1186
rect -3788 1171 -3781 1332
rect -3751 1171 -3743 1328
rect -3684 1320 -3676 1336
rect -3544 1341 -3537 1357
rect -3396 1344 -3389 1360
rect -3544 1333 -3517 1341
rect -3396 1336 -3369 1344
rect -3517 1317 -3509 1333
rect -3738 1302 -3730 1311
rect -3732 1294 -3726 1302
rect -3718 1294 -3668 1302
rect -3646 1298 -3633 1305
rect -3626 1298 -3609 1305
rect -3602 1298 -3587 1305
rect -3571 1299 -3563 1308
rect -3652 1283 -3645 1298
rect -3603 1283 -3596 1298
rect -3562 1291 -3559 1299
rect -3551 1291 -3501 1299
rect -3687 1257 -3648 1263
rect -3630 1259 -3623 1275
rect -3630 1251 -3603 1259
rect -3603 1235 -3595 1251
rect -3657 1218 -3649 1226
rect -3649 1209 -3645 1217
rect -3637 1209 -3617 1217
rect -3609 1209 -3593 1217
rect -3788 1163 -3743 1171
rect -3724 1192 -3710 1198
rect -3703 1192 -3689 1198
rect -3682 1192 -3637 1198
rect -3629 1192 -3619 1198
rect -3610 1192 -3607 1198
rect -3724 1191 -3722 1192
rect -3729 1177 -3722 1191
rect -3680 1177 -3673 1192
rect -3644 1177 -3637 1192
rect -3931 1137 -3925 1144
rect -3881 1142 -3876 1162
rect -3833 1147 -3828 1162
rect -3908 1137 -3876 1142
rect -3908 1125 -3902 1137
rect -3833 1125 -3828 1141
rect -3751 1146 -3743 1163
rect -3707 1153 -3700 1169
rect -3622 1154 -3615 1169
rect -3707 1145 -3680 1153
rect -3680 1129 -3672 1145
rect -3622 1129 -3615 1146
rect -4551 1107 -4354 1110
rect -4366 1102 -4354 1107
rect -4346 1102 -4317 1110
rect -4309 1102 -4275 1110
rect -4266 1102 -4256 1110
rect -4247 1102 -4067 1110
rect -4059 1102 -4031 1110
rect -4023 1102 -3988 1110
rect -3979 1102 -3969 1110
rect -3960 1108 -3940 1110
rect -3928 1108 -3923 1120
rect -3882 1108 -3877 1120
rect -3859 1108 -3853 1120
rect -3734 1111 -3726 1120
rect -3651 1111 -3643 1120
rect -3604 1112 -3595 1209
rect -3436 1146 -3428 1328
rect -3369 1320 -3361 1336
rect -3229 1341 -3222 1357
rect -3229 1333 -3202 1341
rect -3202 1317 -3194 1333
rect -3423 1302 -3415 1311
rect -3417 1294 -3411 1302
rect -3403 1294 -3353 1302
rect -3331 1298 -3318 1305
rect -3311 1298 -3294 1305
rect -3287 1298 -3272 1305
rect -3256 1299 -3248 1308
rect -3337 1283 -3330 1298
rect -3288 1283 -3281 1298
rect -3247 1291 -3244 1299
rect -3236 1291 -3186 1299
rect -3372 1257 -3333 1263
rect -3315 1259 -3308 1275
rect -3315 1251 -3288 1259
rect -3288 1235 -3280 1251
rect -3342 1218 -3334 1226
rect -3334 1209 -3330 1217
rect -3322 1209 -3302 1217
rect -3294 1209 -3278 1217
rect -3409 1192 -3395 1198
rect -3388 1192 -3374 1198
rect -3367 1192 -3322 1198
rect -3314 1192 -3304 1198
rect -3295 1192 -3292 1198
rect -3409 1191 -3407 1192
rect -3414 1177 -3407 1191
rect -3365 1177 -3358 1192
rect -3329 1177 -3322 1192
rect -3392 1153 -3385 1169
rect -3392 1145 -3365 1153
rect -3365 1129 -3357 1145
rect -3307 1129 -3300 1169
rect -3419 1112 -3411 1120
rect -3604 1111 -3411 1112
rect -3336 1111 -3328 1120
rect -3289 1111 -3280 1209
rect -3179 1193 -3174 1380
rect -3267 1187 -3258 1193
rect -3252 1187 -3232 1193
rect -3226 1187 -3205 1193
rect -3199 1187 -3186 1193
rect -3180 1187 -3174 1193
rect -3267 1172 -3262 1187
rect -3194 1172 -3189 1187
rect -3271 1138 -3265 1145
rect -3221 1143 -3216 1163
rect -3173 1147 -3168 1163
rect -3248 1138 -3216 1143
rect -3173 1142 -3155 1147
rect -3248 1126 -3242 1138
rect -3173 1126 -3168 1142
rect -3734 1108 -3722 1111
rect -3960 1102 -3922 1108
rect -3916 1102 -3891 1108
rect -3885 1102 -3869 1108
rect -3863 1102 -3850 1108
rect -3844 1103 -3722 1108
rect -3714 1103 -3685 1111
rect -3677 1103 -3643 1111
rect -3634 1103 -3624 1111
rect -3615 1103 -3407 1111
rect -3399 1103 -3371 1111
rect -3363 1103 -3328 1111
rect -3319 1103 -3309 1111
rect -3300 1109 -3280 1111
rect -3268 1109 -3263 1121
rect -3222 1109 -3217 1121
rect -3199 1109 -3193 1121
rect -3300 1103 -3262 1109
rect -3256 1103 -3231 1109
rect -3225 1103 -3209 1109
rect -3203 1103 -3190 1109
rect -3184 1103 -3176 1109
rect -3844 1102 -3726 1103
rect -4665 1096 -4646 1102
rect -4639 1096 -4619 1102
rect -4612 1096 -4573 1102
rect -4565 1096 -4555 1102
rect -4546 1096 -4541 1102
rect -4665 1081 -4658 1096
rect -4616 1081 -4609 1096
rect -4580 1081 -4573 1096
rect -4488 1086 -4324 1093
rect -4037 1085 -4032 1088
rect -4643 1057 -4636 1073
rect -4643 1049 -4616 1057
rect -4616 1033 -4608 1049
rect -4558 1052 -4551 1073
rect -3692 1070 -3687 1086
rect -3377 1079 -3372 1092
rect -3692 1063 -3188 1070
rect -4558 1044 -4520 1052
rect -4558 1033 -4551 1044
rect -4278 1041 -4265 1048
rect -4258 1041 -4244 1048
rect -4237 1041 -4225 1048
rect -3991 1041 -3978 1048
rect -3971 1041 -3957 1048
rect -3950 1041 -3938 1048
rect -3645 1041 -3632 1048
rect -3625 1041 -3611 1048
rect -3604 1041 -3592 1048
rect -3363 1041 -3350 1048
rect -3343 1041 -3329 1048
rect -3322 1041 -3310 1048
rect -3036 1046 -3023 1053
rect -3016 1046 -3002 1053
rect -2995 1046 -2983 1053
rect -4284 1026 -4277 1041
rect -4235 1026 -4228 1041
rect -4670 1015 -4662 1024
rect -4587 1015 -4579 1024
rect -3997 1026 -3990 1041
rect -3948 1026 -3941 1041
rect -3651 1026 -3644 1041
rect -3602 1026 -3595 1041
rect -3369 1026 -3362 1041
rect -3320 1026 -3313 1041
rect -3042 1031 -3035 1046
rect -2993 1031 -2986 1046
rect -4662 1007 -4658 1015
rect -4650 1007 -4622 1015
rect -4614 1007 -4579 1015
rect -4570 1007 -4560 1015
rect -4551 1007 -4550 1015
rect -4262 1002 -4255 1018
rect -3975 1002 -3968 1018
rect -3629 1002 -3622 1018
rect -3347 1002 -3340 1018
rect -3020 1007 -3013 1023
rect -4348 996 -4285 1001
rect -4665 989 -4646 995
rect -4639 989 -4620 995
rect -4612 989 -4573 995
rect -4565 989 -4555 995
rect -4546 989 -4541 995
rect -4536 989 -4360 995
rect -4262 994 -4235 1002
rect -4215 994 -4190 1002
rect -4061 996 -3998 1001
rect -3975 994 -3948 1002
rect -3928 994 -3903 1002
rect -3715 996 -3652 1001
rect -3629 994 -3602 1002
rect -3582 994 -3557 1002
rect -3433 996 -3370 1001
rect -3347 994 -3320 1002
rect -3300 994 -3275 1002
rect -3106 1001 -3043 1006
rect -3020 999 -2993 1007
rect -2973 999 -2948 1007
rect -4665 974 -4658 989
rect -4616 974 -4609 989
rect -4580 974 -4573 989
rect -4643 950 -4636 966
rect -4558 953 -4551 966
rect -4365 973 -4360 989
rect -4235 978 -4227 994
rect -3948 978 -3940 994
rect -3602 978 -3594 994
rect -3320 978 -3312 994
rect -2993 983 -2985 999
rect -4360 966 -4346 973
rect -4339 966 -4325 973
rect -4318 966 -4304 973
rect -4643 942 -4616 950
rect -4616 926 -4608 942
rect -4558 944 -4496 953
rect -4365 951 -4358 966
rect -4316 951 -4309 966
rect -4289 960 -4281 969
rect -4191 965 -4179 970
rect -4198 963 -4179 965
rect -4172 963 -4158 970
rect -4151 963 -4133 970
rect -4073 966 -4059 973
rect -4052 966 -4038 973
rect -4031 966 -4017 973
rect -4289 952 -4277 960
rect -4269 952 -4224 960
rect -4558 926 -4551 944
rect -4198 948 -4191 963
rect -4149 948 -4142 963
rect -4343 927 -4336 943
rect -4078 951 -4071 966
rect -4029 951 -4022 966
rect -4002 960 -3994 969
rect -3904 965 -3892 970
rect -3911 963 -3892 965
rect -3885 963 -3871 970
rect -3864 966 -3732 970
rect -3727 966 -3713 973
rect -3706 966 -3692 973
rect -3685 966 -3671 973
rect -3864 963 -3725 966
rect -4002 952 -3990 960
rect -3982 952 -3937 960
rect -3911 948 -3904 963
rect -3862 948 -3855 963
rect -4343 919 -4316 927
rect -4670 908 -4662 917
rect -4587 908 -4579 917
rect -4662 900 -4658 908
rect -4650 900 -4622 908
rect -4614 900 -4579 908
rect -4570 900 -4560 908
rect -4551 900 -4550 908
rect -4665 889 -4646 895
rect -4639 889 -4620 895
rect -4612 889 -4573 895
rect -4565 889 -4555 895
rect -4546 889 -4541 895
rect -4665 874 -4658 889
rect -4616 874 -4609 889
rect -4580 874 -4573 889
rect -4681 433 -4675 846
rect -4643 850 -4636 866
rect -4643 842 -4616 850
rect -4616 826 -4608 842
rect -4558 848 -4551 866
rect -4558 841 -4462 848
rect -4558 826 -4551 841
rect -4670 808 -4662 817
rect -4587 808 -4579 817
rect -4662 800 -4658 808
rect -4650 800 -4622 808
rect -4614 800 -4579 808
rect -4570 800 -4560 808
rect -4551 800 -4550 808
rect -4666 774 -4647 780
rect -4640 774 -4623 780
rect -4616 774 -4574 780
rect -4566 774 -4556 780
rect -4547 774 -4541 780
rect -4666 759 -4659 774
rect -4617 759 -4610 774
rect -4581 759 -4574 774
rect -4644 735 -4637 751
rect -4644 727 -4617 735
rect -4617 711 -4609 727
rect -4559 733 -4552 751
rect -4383 747 -4375 911
rect -4316 903 -4308 919
rect -4176 924 -4169 940
rect -4056 927 -4049 943
rect -4176 916 -4149 924
rect -4056 919 -4029 927
rect -4149 900 -4141 916
rect -4370 885 -4362 894
rect -4364 877 -4358 885
rect -4350 877 -4300 885
rect -4278 881 -4265 888
rect -4258 881 -4241 888
rect -4234 881 -4219 888
rect -4203 882 -4195 891
rect -4284 866 -4277 881
rect -4235 866 -4228 881
rect -4194 874 -4191 882
rect -4183 874 -4133 882
rect -4319 840 -4280 846
rect -4262 842 -4255 858
rect -4262 834 -4235 842
rect -4235 818 -4227 834
rect -4289 801 -4281 809
rect -4281 792 -4277 800
rect -4269 792 -4249 800
rect -4241 792 -4225 800
rect -4356 775 -4342 781
rect -4335 775 -4321 781
rect -4314 775 -4269 781
rect -4261 775 -4251 781
rect -4242 775 -4239 781
rect -4356 774 -4354 775
rect -4361 760 -4354 774
rect -4312 760 -4305 775
rect -4276 760 -4269 775
rect -4500 740 -4375 747
rect -4559 726 -4485 733
rect -4383 729 -4375 740
rect -4559 711 -4552 726
rect -4339 736 -4332 752
rect -4254 737 -4247 752
rect -4339 728 -4312 736
rect -4312 712 -4304 728
rect -4254 712 -4247 729
rect -4671 693 -4663 702
rect -4588 693 -4580 702
rect -4366 694 -4358 703
rect -4283 694 -4275 703
rect -4236 695 -4227 792
rect -4096 729 -4088 911
rect -4029 903 -4021 919
rect -3889 924 -3882 940
rect -3889 916 -3862 924
rect -3862 900 -3854 916
rect -4083 885 -4075 894
rect -4077 877 -4071 885
rect -4063 877 -4013 885
rect -3991 881 -3978 888
rect -3971 881 -3954 888
rect -3947 881 -3932 888
rect -3916 882 -3908 891
rect -3997 866 -3990 881
rect -3948 866 -3941 881
rect -3907 874 -3904 882
rect -3896 874 -3846 882
rect -4032 840 -3993 846
rect -3975 842 -3968 858
rect -3975 834 -3948 842
rect -3948 818 -3940 834
rect -4002 801 -3994 809
rect -3994 792 -3990 800
rect -3982 792 -3962 800
rect -3954 792 -3938 800
rect -4069 775 -4055 781
rect -4048 775 -4034 781
rect -4027 775 -3982 781
rect -3974 775 -3964 781
rect -3955 775 -3952 781
rect -4069 774 -4067 775
rect -4074 760 -4067 774
rect -4025 760 -4018 775
rect -3989 760 -3982 775
rect -4052 736 -4045 752
rect -4052 728 -4025 736
rect -4025 712 -4017 728
rect -3967 712 -3960 752
rect -4079 695 -4071 703
rect -4236 694 -4071 695
rect -3996 694 -3988 703
rect -3949 694 -3940 792
rect -3839 776 -3834 963
rect -3732 951 -3725 963
rect -3683 951 -3676 966
rect -3656 960 -3648 969
rect -3558 965 -3546 970
rect -3565 963 -3546 965
rect -3539 963 -3525 970
rect -3518 963 -3500 970
rect -3445 966 -3431 973
rect -3424 966 -3410 973
rect -3403 966 -3389 973
rect -3118 971 -3104 978
rect -3097 971 -3083 978
rect -3076 971 -3062 978
rect -3123 970 -3116 971
rect -3656 952 -3644 960
rect -3636 952 -3591 960
rect -3565 948 -3558 963
rect -3516 948 -3509 963
rect -3710 927 -3703 943
rect -3450 951 -3443 966
rect -3401 951 -3394 966
rect -3374 960 -3366 969
rect -3276 965 -3264 970
rect -3283 963 -3264 965
rect -3257 963 -3243 970
rect -3236 963 -3116 970
rect -3374 952 -3362 960
rect -3354 952 -3309 960
rect -3283 948 -3276 963
rect -3234 948 -3227 963
rect -3710 919 -3683 927
rect -3803 911 -3796 916
rect -3927 770 -3918 776
rect -3912 770 -3892 776
rect -3886 770 -3865 776
rect -3859 770 -3846 776
rect -3840 770 -3834 776
rect -3927 755 -3922 770
rect -3854 755 -3849 770
rect -3931 721 -3925 728
rect -3881 726 -3876 746
rect -3833 730 -3828 746
rect -3908 721 -3876 726
rect -3833 725 -3817 730
rect -3750 729 -3742 911
rect -3683 903 -3675 919
rect -3543 924 -3536 940
rect -3428 927 -3421 943
rect -3543 916 -3516 924
rect -3428 919 -3401 927
rect -3516 900 -3508 916
rect -3737 885 -3729 894
rect -3731 877 -3725 885
rect -3717 877 -3667 885
rect -3645 881 -3632 888
rect -3625 881 -3608 888
rect -3601 881 -3586 888
rect -3570 882 -3562 891
rect -3651 866 -3644 881
rect -3602 866 -3595 881
rect -3561 874 -3558 882
rect -3550 874 -3500 882
rect -3686 840 -3647 846
rect -3629 842 -3622 858
rect -3629 834 -3602 842
rect -3602 818 -3594 834
rect -3656 801 -3648 809
rect -3648 792 -3644 800
rect -3636 792 -3616 800
rect -3608 792 -3592 800
rect -3723 775 -3709 781
rect -3702 775 -3688 781
rect -3681 775 -3636 781
rect -3628 775 -3618 781
rect -3609 775 -3606 781
rect -3723 774 -3721 775
rect -3728 760 -3721 774
rect -3679 760 -3672 775
rect -3643 760 -3636 775
rect -3908 709 -3902 721
rect -3833 709 -3828 725
rect -3796 722 -3750 729
rect -3706 736 -3699 752
rect -3621 737 -3614 752
rect -3706 728 -3679 736
rect -3679 712 -3671 728
rect -3621 712 -3614 729
rect -4366 693 -4354 694
rect -4663 685 -4659 693
rect -4651 685 -4623 693
rect -4615 685 -4580 693
rect -4571 685 -4561 693
rect -4552 686 -4354 693
rect -4346 686 -4317 694
rect -4309 686 -4275 694
rect -4266 686 -4256 694
rect -4247 686 -4067 694
rect -4059 686 -4031 694
rect -4023 686 -3988 694
rect -3979 686 -3969 694
rect -3960 692 -3940 694
rect -3928 692 -3923 704
rect -3882 692 -3877 704
rect -3859 692 -3853 704
rect -3733 694 -3725 703
rect -3650 694 -3642 703
rect -3603 695 -3594 792
rect -3468 729 -3460 911
rect -3401 903 -3393 919
rect -3261 924 -3254 940
rect -3261 916 -3234 924
rect -3234 900 -3226 916
rect -3455 885 -3447 894
rect -3449 877 -3443 885
rect -3435 877 -3385 885
rect -3363 881 -3350 888
rect -3343 881 -3326 888
rect -3319 881 -3304 888
rect -3288 882 -3280 891
rect -3369 866 -3362 881
rect -3320 866 -3313 881
rect -3279 874 -3276 882
rect -3268 874 -3218 882
rect -3404 840 -3365 846
rect -3347 842 -3340 858
rect -3347 834 -3320 842
rect -3320 818 -3312 834
rect -3374 801 -3366 809
rect -3366 792 -3362 800
rect -3354 792 -3334 800
rect -3326 792 -3310 800
rect -3441 775 -3427 781
rect -3420 775 -3406 781
rect -3399 775 -3354 781
rect -3346 775 -3336 781
rect -3327 775 -3324 781
rect -3441 774 -3439 775
rect -3446 760 -3439 774
rect -3397 760 -3390 775
rect -3361 760 -3354 775
rect -3424 736 -3417 752
rect -3424 728 -3397 736
rect -3397 712 -3389 728
rect -3339 712 -3332 752
rect -3451 695 -3443 703
rect -3603 694 -3443 695
rect -3368 694 -3360 703
rect -3321 694 -3312 792
rect -3211 776 -3206 963
rect -3123 956 -3116 963
rect -3074 956 -3067 971
rect -3047 965 -3039 974
rect -2949 970 -2937 975
rect -2956 968 -2937 970
rect -2930 968 -2916 975
rect -2909 968 -2891 975
rect -3047 957 -3035 965
rect -3027 957 -2982 965
rect -2956 953 -2949 968
rect -2907 953 -2900 968
rect -3101 932 -3094 948
rect -3101 924 -3074 932
rect -3169 916 -3141 924
rect -3299 770 -3290 776
rect -3284 770 -3264 776
rect -3258 770 -3237 776
rect -3231 770 -3218 776
rect -3212 770 -3206 776
rect -3299 755 -3294 770
rect -3226 755 -3221 770
rect -3303 721 -3297 728
rect -3253 726 -3248 746
rect -3205 731 -3200 746
rect -3141 734 -3133 916
rect -3074 908 -3066 924
rect -2934 929 -2927 945
rect -2934 921 -2907 929
rect -2907 905 -2899 921
rect -3128 890 -3120 899
rect -3122 882 -3116 890
rect -3108 882 -3058 890
rect -3036 886 -3023 893
rect -3016 886 -2999 893
rect -2992 886 -2977 893
rect -2961 887 -2953 896
rect -3042 871 -3035 886
rect -2993 871 -2986 886
rect -2952 879 -2949 887
rect -2941 879 -2891 887
rect -3077 845 -3038 851
rect -3020 847 -3013 863
rect -3020 839 -2993 847
rect -2993 823 -2985 839
rect -3047 806 -3039 814
rect -3039 797 -3035 805
rect -3027 797 -3007 805
rect -2999 797 -2983 805
rect -3114 780 -3100 786
rect -3093 780 -3079 786
rect -3072 780 -3027 786
rect -3019 780 -3009 786
rect -3000 780 -2997 786
rect -3114 779 -3112 780
rect -3119 765 -3112 779
rect -3070 765 -3063 780
rect -3034 765 -3027 780
rect -3280 721 -3248 726
rect -3205 725 -3188 731
rect -3097 741 -3090 757
rect -3012 741 -3005 757
rect -3097 733 -3070 741
rect -3280 709 -3274 721
rect -3205 709 -3200 725
rect -3070 717 -3062 733
rect -3012 717 -3005 734
rect -3733 692 -3721 694
rect -3960 686 -3922 692
rect -3916 686 -3891 692
rect -3885 686 -3869 692
rect -3863 686 -3850 692
rect -3844 686 -3721 692
rect -3713 686 -3684 694
rect -3676 686 -3642 694
rect -3633 686 -3623 694
rect -3614 686 -3439 694
rect -3431 686 -3403 694
rect -3395 686 -3360 694
rect -3351 686 -3341 694
rect -3332 692 -3312 694
rect -3300 692 -3295 704
rect -3254 692 -3249 704
rect -3231 692 -3225 704
rect -3124 699 -3116 708
rect -3041 699 -3033 708
rect -2994 699 -2985 797
rect -3124 692 -3112 699
rect -3332 686 -3294 692
rect -3288 686 -3263 692
rect -3257 686 -3241 692
rect -3235 686 -3222 692
rect -3216 691 -3112 692
rect -3104 691 -3074 699
rect -3066 691 -3033 699
rect -3024 691 -3014 699
rect -3005 691 -2985 699
rect -3216 686 -3116 691
rect -4552 685 -4551 686
rect -4666 674 -4647 680
rect -4640 674 -4622 680
rect -4614 674 -4574 680
rect -4566 674 -4556 680
rect -4547 674 -4541 680
rect -3077 679 -2841 686
rect -4666 659 -4659 674
rect -4617 659 -4610 674
rect -4581 659 -4574 674
rect -4512 666 -4324 673
rect -4118 663 -4037 671
rect -3691 663 -3686 669
rect -3480 665 -3409 673
rect -4644 635 -4637 651
rect -4644 627 -4617 635
rect -4617 611 -4609 627
rect -4559 634 -4552 651
rect -4559 627 -4473 634
rect -4559 611 -4552 627
rect -4671 593 -4663 602
rect -4588 593 -4580 602
rect -4477 595 -3691 602
rect -4663 585 -4659 593
rect -4651 585 -4623 593
rect -4615 585 -4580 593
rect -4571 585 -4561 593
rect -4552 585 -4551 593
rect -4278 583 -4265 590
rect -4258 583 -4244 590
rect -4237 583 -4225 590
rect -3979 583 -3966 590
rect -3959 583 -3945 590
rect -3938 583 -3926 590
rect -3664 583 -3651 590
rect -3644 583 -3630 590
rect -3623 583 -3611 590
rect -3335 589 -3322 596
rect -3315 589 -3301 596
rect -3294 589 -3282 596
rect -3020 589 -3007 596
rect -3000 589 -2986 596
rect -2979 589 -2967 596
rect -4666 567 -4647 573
rect -4640 567 -4622 573
rect -4615 567 -4574 573
rect -4566 567 -4556 573
rect -4547 567 -4541 573
rect -4284 568 -4277 583
rect -4235 568 -4228 583
rect -4666 552 -4659 567
rect -4617 552 -4610 567
rect -4581 552 -4574 567
rect -3985 568 -3978 583
rect -3936 568 -3929 583
rect -3670 568 -3663 583
rect -3621 568 -3614 583
rect -3341 574 -3334 589
rect -3292 574 -3285 589
rect -3026 574 -3019 589
rect -2977 574 -2970 589
rect -4524 548 -4328 555
rect -4644 528 -4637 544
rect -4644 520 -4617 528
rect -4617 504 -4609 520
rect -4559 524 -4552 544
rect -4262 544 -4255 560
rect -3963 544 -3956 560
rect -3648 544 -3641 560
rect -3319 550 -3312 566
rect -3004 550 -2997 566
rect -3405 544 -3342 549
rect -4351 538 -4285 543
rect -4262 536 -4235 544
rect -4215 536 -4190 544
rect -4052 538 -3986 543
rect -3963 536 -3936 544
rect -3916 536 -3891 544
rect -3734 538 -3671 543
rect -3648 536 -3621 544
rect -3601 536 -3576 544
rect -3319 542 -3292 550
rect -3272 542 -3247 550
rect -3090 544 -3027 549
rect -3004 542 -2932 550
rect -4559 517 -4532 524
rect -4235 520 -4227 536
rect -3936 520 -3928 536
rect -3621 520 -3613 536
rect -3292 526 -3284 542
rect -2977 526 -2969 542
rect -4559 504 -4552 517
rect -4360 508 -4346 515
rect -4339 508 -4322 515
rect -4315 508 -4304 515
rect -4671 486 -4663 495
rect -4588 486 -4580 495
rect -4365 493 -4358 508
rect -4316 493 -4309 508
rect -4289 502 -4281 511
rect -4191 507 -4179 512
rect -4198 505 -4179 507
rect -4172 505 -4158 512
rect -4151 508 -4066 512
rect -4061 508 -4047 515
rect -4040 508 -4026 515
rect -4019 508 -4005 515
rect -4151 505 -4059 508
rect -4289 494 -4277 502
rect -4269 494 -4224 502
rect -4663 478 -4659 486
rect -4651 478 -4623 486
rect -4615 478 -4580 486
rect -4571 478 -4561 486
rect -4552 478 -4551 486
rect -4198 490 -4191 505
rect -4149 490 -4142 505
rect -4666 467 -4647 473
rect -4640 467 -4622 473
rect -4615 467 -4574 473
rect -4566 467 -4556 473
rect -4547 467 -4541 473
rect -4536 467 -4400 473
rect -4343 469 -4336 485
rect -4066 493 -4059 505
rect -4017 493 -4010 508
rect -3990 502 -3982 511
rect -3892 507 -3880 512
rect -3899 505 -3880 507
rect -3873 505 -3859 512
rect -3852 505 -3834 512
rect -3746 508 -3732 515
rect -3725 508 -3711 515
rect -3704 508 -3690 515
rect -3417 514 -3403 521
rect -3396 514 -3382 521
rect -3375 514 -3361 521
rect -3512 512 -3415 514
rect -3990 494 -3978 502
rect -3970 494 -3925 502
rect -3899 490 -3892 505
rect -3850 490 -3843 505
rect -4666 452 -4659 467
rect -4617 452 -4610 467
rect -4581 452 -4574 467
rect -4343 461 -4316 469
rect -4681 21 -4675 427
rect -4644 428 -4637 444
rect -4644 420 -4617 428
rect -4617 404 -4609 420
rect -4559 426 -4552 444
rect -4559 418 -4515 426
rect -4559 404 -4552 418
rect -4671 386 -4663 395
rect -4588 386 -4580 395
rect -4663 378 -4659 386
rect -4651 378 -4623 386
rect -4615 378 -4580 386
rect -4571 378 -4561 386
rect -4552 378 -4551 386
rect -4666 364 -4647 370
rect -4640 364 -4624 370
rect -4617 364 -4574 370
rect -4566 364 -4556 370
rect -4547 364 -4541 370
rect -4666 349 -4659 364
rect -4617 349 -4610 364
rect -4581 349 -4574 364
rect -4644 325 -4637 341
rect -4559 327 -4552 341
rect -4644 317 -4617 325
rect -4617 301 -4609 317
rect -4559 319 -4429 327
rect -4559 301 -4552 319
rect -4383 304 -4375 453
rect -4316 445 -4308 461
rect -4176 466 -4169 482
rect -4044 469 -4037 485
rect -3751 493 -3744 508
rect -3702 493 -3695 508
rect -3675 502 -3667 511
rect -3577 507 -3565 512
rect -3584 505 -3565 507
rect -3558 505 -3544 512
rect -3537 507 -3415 512
rect -3537 505 -3507 507
rect -3675 494 -3663 502
rect -3655 494 -3610 502
rect -3584 490 -3577 505
rect -3535 490 -3528 505
rect -4176 458 -4149 466
rect -4149 442 -4141 458
rect -4370 427 -4362 436
rect -4044 461 -4017 469
rect -4364 419 -4358 427
rect -4350 419 -4300 427
rect -4278 423 -4265 430
rect -4258 423 -4241 430
rect -4234 423 -4219 430
rect -4203 424 -4195 433
rect -4284 408 -4277 423
rect -4235 408 -4228 423
rect -4194 416 -4191 424
rect -4183 416 -4133 424
rect -4319 382 -4280 388
rect -4262 384 -4255 400
rect -4262 376 -4235 384
rect -4235 360 -4227 376
rect -4289 343 -4281 351
rect -4281 334 -4277 342
rect -4269 334 -4249 342
rect -4241 334 -4225 342
rect -4489 298 -4375 304
rect -4671 283 -4663 292
rect -4588 283 -4580 292
rect -4663 275 -4659 283
rect -4651 275 -4623 283
rect -4615 275 -4580 283
rect -4571 275 -4561 283
rect -4552 275 -4399 283
rect -4666 264 -4647 270
rect -4640 264 -4622 270
rect -4615 264 -4574 270
rect -4566 264 -4556 270
rect -4547 264 -4541 270
rect -4666 249 -4659 264
rect -4617 249 -4610 264
rect -4581 249 -4574 264
rect -4644 225 -4637 241
rect -4644 217 -4617 225
rect -4617 201 -4609 217
rect -4559 215 -4552 241
rect -4406 236 -4399 275
rect -4383 271 -4375 298
rect -4356 317 -4342 323
rect -4335 317 -4321 323
rect -4314 317 -4269 323
rect -4261 317 -4251 323
rect -4242 317 -4239 323
rect -4356 316 -4354 317
rect -4361 302 -4354 316
rect -4312 302 -4305 317
rect -4276 302 -4269 317
rect -4339 278 -4332 294
rect -4254 279 -4247 294
rect -4339 270 -4312 278
rect -4312 254 -4304 270
rect -4254 254 -4247 271
rect -4366 236 -4358 245
rect -4283 236 -4275 245
rect -4236 237 -4227 334
rect -4216 271 -4126 279
rect -4084 271 -4076 458
rect -4017 445 -4009 461
rect -3877 466 -3870 482
rect -3729 469 -3722 485
rect -3877 458 -3850 466
rect -3729 461 -3702 469
rect -3850 442 -3842 458
rect -4071 427 -4063 436
rect -4065 419 -4059 427
rect -4051 419 -4001 427
rect -3979 423 -3966 430
rect -3959 423 -3942 430
rect -3935 423 -3920 430
rect -3904 424 -3896 433
rect -3985 408 -3978 423
rect -3936 408 -3929 423
rect -3895 416 -3892 424
rect -3884 416 -3834 424
rect -4020 382 -3981 388
rect -3963 384 -3956 400
rect -3963 376 -3936 384
rect -3936 360 -3928 376
rect -3990 343 -3982 351
rect -3982 334 -3978 342
rect -3970 334 -3950 342
rect -3942 334 -3926 342
rect -4057 317 -4043 323
rect -4036 317 -4022 323
rect -4015 317 -3970 323
rect -3962 317 -3952 323
rect -3943 317 -3940 323
rect -4057 316 -4055 317
rect -4062 302 -4055 316
rect -4013 302 -4006 317
rect -3977 302 -3970 317
rect -4040 278 -4033 294
rect -3955 279 -3948 294
rect -4040 270 -4013 278
rect -4013 254 -4005 270
rect -3955 254 -3948 271
rect -4067 237 -4059 245
rect -4236 236 -4059 237
rect -3984 236 -3976 245
rect -3937 237 -3928 334
rect -3769 271 -3761 453
rect -3702 445 -3694 461
rect -3562 466 -3555 482
rect -3562 458 -3535 466
rect -3535 442 -3527 458
rect -3756 427 -3748 436
rect -3750 419 -3744 427
rect -3736 419 -3686 427
rect -3664 423 -3651 430
rect -3644 423 -3627 430
rect -3620 423 -3605 430
rect -3589 424 -3581 433
rect -3670 408 -3663 423
rect -3621 408 -3614 423
rect -3580 416 -3577 424
rect -3569 416 -3519 424
rect -3705 382 -3666 388
rect -3648 384 -3641 400
rect -3648 376 -3621 384
rect -3621 360 -3613 376
rect -3675 343 -3667 351
rect -3667 334 -3663 342
rect -3655 334 -3635 342
rect -3627 334 -3611 342
rect -3742 317 -3728 323
rect -3721 317 -3707 323
rect -3700 317 -3655 323
rect -3647 317 -3637 323
rect -3628 317 -3625 323
rect -3742 316 -3740 317
rect -3747 302 -3740 316
rect -3698 302 -3691 317
rect -3662 302 -3655 317
rect -3725 278 -3718 294
rect -3725 270 -3698 278
rect -3698 254 -3690 270
rect -3640 254 -3633 294
rect -3752 237 -3744 245
rect -3937 236 -3744 237
rect -3669 236 -3661 245
rect -3622 236 -3613 334
rect -3512 298 -3507 505
rect -3422 499 -3415 507
rect -3373 499 -3366 514
rect -3346 508 -3338 517
rect -3248 513 -3236 518
rect -3255 511 -3236 513
rect -3229 511 -3215 518
rect -3208 511 -3190 518
rect -3102 514 -3088 521
rect -3081 514 -3067 521
rect -3060 514 -3046 521
rect -3346 500 -3334 508
rect -3326 500 -3281 508
rect -3255 496 -3248 511
rect -3206 496 -3199 511
rect -3400 475 -3393 491
rect -3107 499 -3100 514
rect -3058 499 -3051 514
rect -3031 508 -3023 517
rect -2933 513 -2921 518
rect -2940 511 -2921 513
rect -2914 511 -2900 518
rect -2893 511 -2863 518
rect -3031 500 -3019 508
rect -3011 500 -2966 508
rect -2940 496 -2933 511
rect -2891 496 -2884 511
rect -3400 467 -3373 475
rect -3600 292 -3591 298
rect -3585 292 -3565 298
rect -3559 292 -3538 298
rect -3532 292 -3519 298
rect -3513 292 -3507 298
rect -3600 277 -3595 292
rect -3527 277 -3522 292
rect -3468 277 -3460 458
rect -3440 277 -3432 459
rect -3373 451 -3365 467
rect -3233 472 -3226 488
rect -3085 475 -3078 491
rect -3233 464 -3206 472
rect -3085 467 -3058 475
rect -3206 448 -3198 464
rect -3427 433 -3419 442
rect -3421 425 -3415 433
rect -3407 425 -3357 433
rect -3335 429 -3322 436
rect -3315 429 -3298 436
rect -3291 429 -3276 436
rect -3260 430 -3252 439
rect -3341 414 -3334 429
rect -3292 414 -3285 429
rect -3251 422 -3248 430
rect -3240 422 -3190 430
rect -3376 388 -3337 394
rect -3319 390 -3312 406
rect -3319 382 -3292 390
rect -3292 366 -3284 382
rect -3346 349 -3338 357
rect -3338 340 -3334 348
rect -3326 340 -3306 348
rect -3298 340 -3282 348
rect -3413 323 -3399 329
rect -3392 323 -3378 329
rect -3371 323 -3326 329
rect -3318 323 -3308 329
rect -3299 323 -3296 329
rect -3413 322 -3411 323
rect -3418 308 -3411 322
rect -3369 308 -3362 323
rect -3333 308 -3326 323
rect -3468 270 -3440 277
rect -3396 284 -3389 300
rect -3311 285 -3304 300
rect -3396 276 -3369 284
rect -3604 243 -3598 250
rect -3554 248 -3549 268
rect -3506 253 -3501 268
rect -3369 260 -3361 276
rect -3311 260 -3304 277
rect -3581 243 -3549 248
rect -3506 246 -3488 253
rect -4406 228 -4354 236
rect -4346 228 -4326 236
rect -4318 228 -4275 236
rect -4266 228 -4256 236
rect -4247 228 -4055 236
rect -4047 228 -4018 236
rect -4010 228 -3976 236
rect -3967 228 -3957 236
rect -3948 228 -3740 236
rect -3732 228 -3703 236
rect -3695 228 -3661 236
rect -3652 228 -3642 236
rect -3633 228 -3613 236
rect -3581 231 -3575 243
rect -3506 231 -3501 246
rect -4466 219 -4025 225
rect -4559 208 -4484 215
rect -4278 209 -4265 216
rect -4258 209 -4244 216
rect -4237 209 -4225 216
rect -3620 214 -3613 228
rect -3601 214 -3596 226
rect -3555 214 -3550 226
rect -3423 242 -3415 251
rect -3340 242 -3332 251
rect -3293 243 -3284 340
rect -3125 277 -3117 459
rect -3058 451 -3050 467
rect -2918 472 -2911 488
rect -2918 464 -2891 472
rect -2891 448 -2883 464
rect -3112 433 -3104 442
rect -3106 425 -3100 433
rect -3092 425 -3042 433
rect -3020 429 -3007 436
rect -3000 429 -2983 436
rect -2976 429 -2961 436
rect -2945 430 -2937 439
rect -3026 414 -3019 429
rect -2977 414 -2970 429
rect -2936 422 -2933 430
rect -2925 422 -2875 430
rect -3061 388 -3022 394
rect -3004 390 -2997 406
rect -3004 382 -2977 390
rect -2977 366 -2969 382
rect -3031 349 -3023 357
rect -3023 340 -3019 348
rect -3011 340 -2991 348
rect -2983 340 -2967 348
rect -3098 323 -3084 329
rect -3077 323 -3063 329
rect -3056 323 -3011 329
rect -3003 323 -2993 329
rect -2984 323 -2981 329
rect -3098 322 -3096 323
rect -3103 308 -3096 322
rect -3054 308 -3047 323
rect -3018 308 -3011 323
rect -3081 284 -3074 300
rect -3081 276 -3054 284
rect -3054 260 -3046 276
rect -2996 260 -2989 300
rect -3108 243 -3100 251
rect -3293 242 -3100 243
rect -3025 242 -3017 251
rect -2978 242 -2969 340
rect -2868 304 -2863 511
rect -2956 298 -2947 304
rect -2941 298 -2921 304
rect -2915 298 -2894 304
rect -2888 298 -2875 304
rect -2869 298 -2863 304
rect -2956 283 -2951 298
rect -2883 283 -2878 298
rect -2960 249 -2954 256
rect -2910 254 -2905 274
rect -2862 260 -2857 274
rect -2848 260 -2841 679
rect -2937 249 -2905 254
rect -2862 253 -2841 260
rect -3423 234 -3411 242
rect -3403 234 -3374 242
rect -3366 234 -3332 242
rect -3323 234 -3313 242
rect -3304 234 -3096 242
rect -3088 234 -3060 242
rect -3052 234 -3017 242
rect -3008 234 -2998 242
rect -2989 234 -2969 242
rect -2937 237 -2931 249
rect -2862 237 -2857 253
rect -3532 214 -3526 226
rect -3423 214 -3415 234
rect -4559 201 -4552 208
rect -4284 194 -4277 209
rect -4235 194 -4228 209
rect -3620 208 -3595 214
rect -3589 208 -3564 214
rect -3558 208 -3542 214
rect -3536 208 -3523 214
rect -3517 208 -3415 214
rect -4084 199 -3710 207
rect -3381 196 -3376 217
rect -2976 220 -2969 234
rect -2957 220 -2952 232
rect -2911 220 -2906 232
rect -2888 220 -2882 232
rect -2976 214 -2951 220
rect -2945 214 -2920 220
rect -2914 214 -2898 220
rect -2892 214 -2879 220
rect -2873 214 -2865 220
rect -4671 183 -4663 192
rect -4588 183 -4580 192
rect -4119 187 -3376 196
rect -3256 206 -3066 211
rect -4663 175 -4659 183
rect -4651 175 -4623 183
rect -4615 175 -4580 183
rect -4571 175 -4561 183
rect -4552 175 -4551 183
rect -4524 172 -4328 178
rect -4262 170 -4255 186
rect -3947 176 -3934 183
rect -3927 176 -3913 183
rect -3906 176 -3894 183
rect -3632 176 -3619 183
rect -3612 176 -3598 183
rect -3591 176 -3579 183
rect -4348 164 -4285 169
rect -4666 157 -4647 163
rect -4640 157 -4622 163
rect -4615 157 -4574 163
rect -4566 157 -4556 163
rect -4547 157 -4541 163
rect -4536 157 -4360 163
rect -4262 162 -4235 170
rect -4215 162 -4190 170
rect -4666 142 -4659 157
rect -4617 142 -4610 157
rect -4581 142 -4574 157
rect -4644 118 -4637 134
rect -4644 110 -4617 118
rect -4617 94 -4609 110
rect -4559 116 -4552 134
rect -4365 141 -4360 157
rect -4235 146 -4227 162
rect -3953 161 -3946 176
rect -3904 161 -3897 176
rect -3638 161 -3631 176
rect -3589 161 -3582 176
rect -4360 134 -4346 141
rect -4339 134 -4321 141
rect -4314 134 -4304 141
rect -4365 119 -4358 134
rect -4316 119 -4309 134
rect -4289 128 -4281 137
rect -4191 133 -4179 138
rect -4198 131 -4179 133
rect -4172 131 -4158 138
rect -4151 131 -4029 138
rect -3931 137 -3924 153
rect -3616 137 -3609 153
rect -4017 131 -3954 136
rect -4289 120 -4277 128
rect -4269 120 -4224 128
rect -4559 109 -4501 116
rect -4198 116 -4191 131
rect -4149 116 -4142 131
rect -4559 94 -4552 109
rect -4343 95 -4336 111
rect -4034 108 -4029 131
rect -3931 129 -3904 137
rect -3884 129 -3859 137
rect -3702 131 -3639 136
rect -3616 129 -3589 137
rect -3569 129 -3544 137
rect -3904 113 -3896 129
rect -3589 113 -3581 129
rect -4343 87 -4316 95
rect -4671 76 -4663 85
rect -4588 76 -4580 85
rect -4455 79 -4383 86
rect -4663 68 -4659 76
rect -4651 68 -4623 76
rect -4615 68 -4580 76
rect -4571 68 -4561 76
rect -4552 68 -4551 76
rect -4666 57 -4647 63
rect -4640 57 -4623 63
rect -4616 57 -4574 63
rect -4566 57 -4556 63
rect -4547 57 -4541 63
rect -4666 42 -4659 57
rect -4617 42 -4610 57
rect -4581 42 -4574 57
rect -4644 18 -4637 34
rect -4644 10 -4617 18
rect -4617 -6 -4609 10
rect -4559 -6 -4552 34
rect -4671 -24 -4663 -15
rect -4588 -24 -4580 -15
rect -4663 -32 -4659 -24
rect -4651 -32 -4623 -24
rect -4615 -32 -4580 -24
rect -4571 -32 -4561 -24
rect -4552 -32 -4551 -24
rect -4562 -137 -4551 -32
rect -4383 -103 -4375 79
rect -4316 71 -4308 87
rect -4176 92 -4169 108
rect -4029 101 -4015 108
rect -4008 101 -3994 108
rect -3987 101 -3973 108
rect -4176 84 -4149 92
rect -4141 84 -4127 92
rect -4119 84 -4072 92
rect -4034 86 -4027 101
rect -3985 86 -3978 101
rect -3958 95 -3950 104
rect -3860 100 -3848 105
rect -3867 98 -3848 100
rect -3841 98 -3827 105
rect -3820 98 -3802 105
rect -3714 101 -3700 108
rect -3693 101 -3679 108
rect -3672 101 -3658 108
rect -3958 87 -3946 95
rect -3938 87 -3893 95
rect -4149 68 -4141 84
rect -3867 83 -3860 98
rect -3818 83 -3811 98
rect -4370 53 -4362 62
rect -4012 62 -4005 78
rect -3719 86 -3712 101
rect -3670 86 -3663 101
rect -3643 95 -3635 104
rect -3545 100 -3533 105
rect -3552 98 -3533 100
rect -3526 98 -3512 105
rect -3505 98 -3475 105
rect -3643 87 -3631 95
rect -3623 87 -3578 95
rect -3552 83 -3545 98
rect -3503 83 -3496 98
rect -4364 45 -4358 53
rect -4350 45 -4300 53
rect -4278 49 -4265 56
rect -4258 49 -4241 56
rect -4234 49 -4219 56
rect -4203 50 -4195 59
rect -4012 54 -3985 62
rect -4284 34 -4277 49
rect -4235 34 -4228 49
rect -4194 42 -4191 50
rect -4183 42 -4133 50
rect -4319 8 -4280 14
rect -4262 10 -4255 26
rect -4262 2 -4235 10
rect -4235 -14 -4227 2
rect -4289 -31 -4281 -23
rect -4281 -40 -4277 -32
rect -4269 -40 -4249 -32
rect -4241 -40 -4225 -32
rect -4356 -57 -4342 -51
rect -4335 -57 -4321 -51
rect -4314 -57 -4269 -51
rect -4261 -57 -4251 -51
rect -4242 -57 -4239 -51
rect -4356 -58 -4354 -57
rect -4361 -72 -4354 -58
rect -4312 -72 -4305 -57
rect -4276 -72 -4269 -57
rect -4339 -96 -4332 -80
rect -4254 -95 -4247 -80
rect -4339 -104 -4312 -96
rect -4312 -120 -4304 -104
rect -4254 -120 -4247 -103
rect -4366 -137 -4358 -129
rect -4562 -138 -4358 -137
rect -4283 -138 -4275 -129
rect -4236 -136 -4227 -40
rect -4216 -103 -4092 -95
rect -4052 -136 -4044 46
rect -3985 38 -3977 54
rect -3845 59 -3838 75
rect -3697 62 -3690 78
rect -3845 51 -3818 59
rect -3697 54 -3670 62
rect -3818 35 -3810 51
rect -4039 20 -4031 29
rect -4033 12 -4027 20
rect -4019 12 -3969 20
rect -3947 16 -3934 23
rect -3927 16 -3910 23
rect -3903 16 -3888 23
rect -3872 17 -3864 26
rect -3953 1 -3946 16
rect -3904 1 -3897 16
rect -3863 9 -3860 17
rect -3852 9 -3802 17
rect -3988 -25 -3949 -19
rect -3931 -23 -3924 -7
rect -3931 -31 -3904 -23
rect -3904 -47 -3896 -31
rect -3958 -64 -3950 -56
rect -3950 -73 -3946 -65
rect -3938 -73 -3918 -65
rect -3910 -73 -3894 -65
rect -4025 -90 -4011 -84
rect -4004 -90 -3990 -84
rect -3983 -90 -3938 -84
rect -3930 -90 -3920 -84
rect -3911 -90 -3908 -84
rect -4025 -91 -4023 -90
rect -4030 -105 -4023 -91
rect -3981 -105 -3974 -90
rect -3945 -105 -3938 -90
rect -4236 -138 -4077 -136
rect -4562 -146 -4354 -138
rect -4346 -146 -4326 -138
rect -4318 -146 -4275 -138
rect -4266 -146 -4256 -138
rect -4247 -146 -4077 -138
rect -4066 -143 -4052 -136
rect -4008 -129 -4001 -113
rect -3923 -128 -3916 -113
rect -4008 -137 -3981 -129
rect -4562 -511 -4552 -146
rect -4477 -157 -4093 -149
rect -4278 -167 -4265 -160
rect -4258 -167 -4244 -160
rect -4237 -167 -4225 -160
rect -4284 -182 -4277 -167
rect -4235 -182 -4228 -167
rect -4494 -199 -4328 -194
rect -4262 -206 -4255 -190
rect -4101 -192 -4093 -157
rect -4085 -171 -4077 -146
rect -3981 -153 -3973 -137
rect -3923 -153 -3916 -136
rect -4035 -171 -4027 -162
rect -3952 -171 -3944 -162
rect -3905 -170 -3896 -73
rect -3737 -136 -3729 46
rect -3670 38 -3662 54
rect -3530 59 -3523 75
rect -3530 51 -3503 59
rect -3503 35 -3495 51
rect -3724 20 -3716 29
rect -3718 12 -3712 20
rect -3704 12 -3654 20
rect -3632 16 -3619 23
rect -3612 16 -3595 23
rect -3588 16 -3573 23
rect -3557 17 -3549 26
rect -3638 1 -3631 16
rect -3589 1 -3582 16
rect -3548 9 -3545 17
rect -3537 9 -3487 17
rect -3673 -25 -3634 -19
rect -3616 -23 -3609 -7
rect -3616 -31 -3589 -23
rect -3589 -47 -3581 -31
rect -3643 -64 -3635 -56
rect -3635 -73 -3631 -65
rect -3623 -73 -3603 -65
rect -3595 -73 -3579 -65
rect -3710 -90 -3696 -84
rect -3689 -90 -3675 -84
rect -3668 -90 -3623 -84
rect -3615 -90 -3605 -84
rect -3596 -90 -3593 -84
rect -3710 -91 -3708 -90
rect -3715 -105 -3708 -91
rect -3666 -105 -3659 -90
rect -3630 -105 -3623 -90
rect -3693 -129 -3686 -113
rect -3693 -137 -3666 -129
rect -3666 -153 -3658 -137
rect -3608 -153 -3601 -113
rect -3720 -170 -3712 -162
rect -3905 -171 -3712 -170
rect -3637 -171 -3629 -162
rect -3590 -171 -3581 -73
rect -3480 -109 -3475 98
rect -3568 -115 -3559 -109
rect -3553 -115 -3533 -109
rect -3527 -115 -3506 -109
rect -3500 -115 -3487 -109
rect -3481 -115 -3475 -109
rect -3568 -130 -3563 -115
rect -3495 -130 -3490 -115
rect -3572 -164 -3566 -157
rect -3522 -159 -3517 -139
rect -3474 -154 -3469 -139
rect -3256 -154 -3250 206
rect -3549 -164 -3517 -159
rect -3474 -160 -3250 -154
rect -4085 -179 -4023 -171
rect -4015 -179 -3986 -171
rect -3978 -179 -3944 -171
rect -3935 -179 -3925 -171
rect -3916 -179 -3708 -171
rect -3700 -179 -3672 -171
rect -3664 -179 -3629 -171
rect -3620 -179 -3610 -171
rect -3601 -179 -3581 -171
rect -3549 -176 -3543 -164
rect -3474 -176 -3469 -160
rect -4101 -199 -3993 -192
rect -3588 -193 -3581 -179
rect -3569 -193 -3564 -181
rect -3523 -193 -3518 -181
rect -3500 -193 -3494 -181
rect -3588 -199 -3563 -193
rect -3557 -199 -3532 -193
rect -3526 -199 -3510 -193
rect -3504 -199 -3491 -193
rect -3485 -199 -3477 -193
rect -4348 -212 -4285 -207
rect -4262 -214 -4235 -206
rect -4215 -214 -4190 -206
rect -3678 -209 -3673 -205
rect -4235 -230 -4227 -214
rect -4536 -242 -4365 -235
rect -4360 -242 -4346 -235
rect -4339 -242 -4321 -235
rect -4314 -242 -4304 -235
rect -4365 -257 -4358 -242
rect -4316 -257 -4309 -242
rect -4289 -248 -4281 -239
rect -4191 -243 -4179 -238
rect -4198 -245 -4179 -243
rect -4172 -245 -4158 -238
rect -4151 -245 -4133 -238
rect -4289 -256 -4277 -248
rect -4269 -256 -4224 -248
rect -4198 -260 -4191 -245
rect -4149 -260 -4142 -245
rect -4343 -281 -4336 -265
rect -4343 -289 -4316 -281
rect -4507 -297 -4383 -290
rect -4383 -479 -4375 -297
rect -4316 -305 -4308 -289
rect -4176 -284 -4169 -268
rect -4176 -292 -4149 -284
rect -4149 -308 -4141 -292
rect -4370 -323 -4362 -314
rect -4364 -331 -4358 -323
rect -4350 -331 -4300 -323
rect -4278 -327 -4265 -320
rect -4258 -327 -4241 -320
rect -4234 -327 -4219 -320
rect -4203 -326 -4195 -317
rect -4284 -342 -4277 -327
rect -4235 -342 -4228 -327
rect -4194 -334 -4191 -326
rect -4183 -334 -4133 -326
rect -4319 -368 -4280 -362
rect -4262 -366 -4255 -350
rect -4262 -374 -4235 -366
rect -4235 -390 -4227 -374
rect -4289 -407 -4281 -399
rect -4281 -416 -4277 -408
rect -4269 -416 -4249 -408
rect -4241 -416 -4225 -408
rect -4356 -433 -4342 -427
rect -4335 -433 -4321 -427
rect -4314 -433 -4269 -427
rect -4261 -433 -4251 -427
rect -4242 -433 -4239 -427
rect -4356 -434 -4354 -433
rect -4361 -448 -4354 -434
rect -4312 -448 -4305 -433
rect -4276 -448 -4269 -433
rect -4339 -472 -4332 -456
rect -4254 -471 -4247 -456
rect -4339 -480 -4312 -472
rect -4312 -496 -4304 -480
rect -4254 -496 -4247 -479
rect -4366 -511 -4358 -505
rect -4562 -514 -4358 -511
rect -4283 -514 -4275 -505
rect -4236 -514 -4227 -416
rect -4562 -517 -4354 -514
rect -4563 -522 -4354 -517
rect -4346 -522 -4326 -514
rect -4318 -522 -4275 -514
rect -4266 -522 -4256 -514
rect -4247 -522 -4227 -514
<< m2contact >>
rect -4541 1606 -4536 1612
rect -4670 1517 -4662 1525
rect -4431 1522 -4425 1528
rect -4541 1506 -4536 1512
rect -4496 1457 -4488 1465
rect -4284 1457 -4278 1464
rect -4225 1457 -4219 1464
rect -3997 1457 -3991 1464
rect -3938 1457 -3932 1464
rect -3652 1458 -3646 1465
rect -3593 1458 -3587 1465
rect -3337 1458 -3331 1465
rect -3278 1458 -3272 1465
rect -4670 1417 -4662 1425
rect -4541 1399 -4536 1405
rect -4365 1382 -4360 1389
rect -4304 1382 -4298 1389
rect -4198 1381 -4191 1386
rect -4078 1382 -4073 1389
rect -4017 1382 -4011 1389
rect -4224 1368 -4219 1376
rect -4508 1350 -4500 1358
rect -3911 1381 -3904 1386
rect -3733 1383 -3728 1390
rect -3672 1383 -3666 1390
rect -3937 1368 -3932 1376
rect -4670 1310 -4662 1318
rect -4541 1299 -4536 1305
rect -4530 1250 -4524 1257
rect -4670 1210 -4662 1218
rect -4541 1196 -4536 1202
rect -4370 1293 -4364 1301
rect -4284 1297 -4278 1304
rect -4203 1290 -4194 1298
rect -4289 1208 -4281 1217
rect -4225 1208 -4219 1216
rect -4361 1190 -4356 1197
rect -4254 1145 -4247 1153
rect -4670 1107 -4662 1115
rect -4083 1293 -4077 1301
rect -3997 1297 -3991 1304
rect -3916 1290 -3907 1298
rect -4002 1208 -3994 1217
rect -3938 1208 -3932 1216
rect -4074 1190 -4069 1197
rect -3566 1382 -3559 1387
rect -3418 1383 -3413 1390
rect -3357 1383 -3351 1390
rect -3592 1369 -3587 1377
rect -3251 1382 -3244 1387
rect -3277 1369 -3272 1377
rect -3738 1294 -3732 1302
rect -3652 1298 -3646 1305
rect -3571 1291 -3562 1299
rect -3657 1209 -3649 1218
rect -3593 1209 -3587 1217
rect -3729 1191 -3724 1198
rect -3937 1137 -3931 1144
rect -3833 1141 -3828 1147
rect -3622 1146 -3615 1154
rect -3423 1294 -3417 1302
rect -3337 1298 -3331 1305
rect -3256 1291 -3247 1299
rect -3342 1209 -3334 1218
rect -3278 1209 -3272 1217
rect -3414 1191 -3409 1198
rect -3277 1138 -3271 1145
rect -3155 1142 -3149 1147
rect -4541 1096 -4536 1102
rect -4496 1086 -4488 1093
rect -4037 1080 -4032 1085
rect -3377 1073 -3372 1079
rect -3188 1063 -3181 1070
rect -4520 1044 -4512 1052
rect -4284 1041 -4278 1048
rect -4225 1041 -4219 1048
rect -3997 1041 -3991 1048
rect -3938 1041 -3932 1048
rect -3651 1041 -3645 1048
rect -3592 1041 -3586 1048
rect -3369 1041 -3363 1048
rect -3310 1041 -3304 1048
rect -3042 1046 -3036 1053
rect -2983 1046 -2977 1053
rect -4670 1007 -4662 1015
rect -4541 989 -4536 995
rect -4365 966 -4360 973
rect -4304 966 -4298 973
rect -4496 944 -4489 953
rect -4198 965 -4191 970
rect -4078 966 -4073 973
rect -4017 966 -4011 973
rect -4224 952 -4219 960
rect -3911 965 -3904 970
rect -3732 966 -3727 973
rect -3671 966 -3665 973
rect -3937 952 -3932 960
rect -4670 900 -4662 908
rect -4541 889 -4536 895
rect -4462 841 -4455 848
rect -4670 800 -4662 808
rect -4541 774 -4536 780
rect -4370 877 -4364 885
rect -4284 881 -4278 888
rect -4203 874 -4194 882
rect -4289 792 -4281 801
rect -4225 792 -4219 800
rect -4361 774 -4356 781
rect -4508 740 -4500 747
rect -4485 726 -4477 733
rect -4254 729 -4247 737
rect -4083 877 -4077 885
rect -3997 881 -3991 888
rect -3916 874 -3907 882
rect -4002 792 -3994 801
rect -3938 792 -3932 800
rect -4074 774 -4069 781
rect -3565 965 -3558 970
rect -3450 966 -3445 973
rect -3389 966 -3383 973
rect -3123 971 -3118 978
rect -3062 971 -3056 978
rect -3591 952 -3586 960
rect -3283 965 -3276 970
rect -3309 952 -3304 960
rect -3803 905 -3796 911
rect -3937 721 -3931 728
rect -3817 725 -3811 730
rect -3737 877 -3731 885
rect -3651 881 -3645 888
rect -3570 874 -3561 882
rect -3656 792 -3648 801
rect -3592 792 -3586 800
rect -3728 774 -3723 781
rect -3803 722 -3796 729
rect -3621 729 -3614 737
rect -4671 685 -4663 693
rect -3455 877 -3449 885
rect -3369 881 -3363 888
rect -3288 874 -3279 882
rect -3374 792 -3366 801
rect -3310 792 -3304 800
rect -3446 774 -3441 781
rect -2956 970 -2949 975
rect -2982 957 -2977 965
rect -3309 721 -3303 728
rect -3128 882 -3122 890
rect -3042 886 -3036 893
rect -2961 879 -2952 887
rect -3047 797 -3039 806
rect -2983 797 -2977 805
rect -3119 779 -3114 786
rect -3188 725 -3181 731
rect -3012 734 -3005 741
rect -4541 674 -4536 680
rect -4520 666 -4512 673
rect -4126 663 -4118 671
rect -3488 665 -3480 673
rect -3691 657 -3686 663
rect -4473 627 -4466 634
rect -4485 595 -4477 602
rect -3691 595 -3686 602
rect -4671 585 -4663 593
rect -4284 583 -4278 590
rect -4225 583 -4219 590
rect -3985 583 -3979 590
rect -3926 583 -3920 590
rect -3670 583 -3664 590
rect -3611 583 -3605 590
rect -3341 589 -3335 596
rect -3282 589 -3276 596
rect -3026 589 -3020 596
rect -2967 589 -2961 596
rect -4541 567 -4536 573
rect -4530 548 -4524 555
rect -4532 517 -4524 524
rect -4365 508 -4360 515
rect -4304 508 -4298 515
rect -4198 507 -4191 512
rect -4066 508 -4061 515
rect -4005 508 -3999 515
rect -4224 494 -4219 502
rect -4671 478 -4663 486
rect -4541 467 -4536 473
rect -4400 467 -4395 473
rect -3899 507 -3892 512
rect -3751 508 -3746 515
rect -3690 508 -3684 515
rect -3422 514 -3417 521
rect -3361 514 -3355 521
rect -3925 494 -3920 502
rect -4515 418 -4507 426
rect -4671 378 -4663 386
rect -4541 364 -4536 370
rect -4429 319 -4421 327
rect -3584 507 -3577 512
rect -3610 494 -3605 502
rect -4370 419 -4364 427
rect -4284 423 -4278 430
rect -4203 416 -4194 424
rect -4289 334 -4281 343
rect -4225 334 -4219 342
rect -4496 298 -4489 304
rect -4671 275 -4663 283
rect -4541 264 -4536 270
rect -4361 316 -4356 323
rect -4254 271 -4247 279
rect -4223 271 -4216 279
rect -4126 271 -4118 279
rect -4071 419 -4065 427
rect -3985 423 -3979 430
rect -3904 416 -3895 424
rect -3990 334 -3982 343
rect -3926 334 -3920 342
rect -4062 316 -4057 323
rect -3955 271 -3948 279
rect -3756 419 -3750 427
rect -3670 423 -3664 430
rect -3589 416 -3580 424
rect -3675 334 -3667 343
rect -3611 334 -3605 342
rect -3747 316 -3742 323
rect -3255 513 -3248 518
rect -3107 514 -3102 521
rect -3046 514 -3040 521
rect -3281 500 -3276 508
rect -2940 513 -2933 518
rect -2966 500 -2961 508
rect -3427 425 -3421 433
rect -3341 429 -3335 436
rect -3260 422 -3251 430
rect -3346 340 -3338 349
rect -3282 340 -3276 348
rect -3418 322 -3413 329
rect -3610 243 -3604 250
rect -3311 277 -3304 285
rect -3488 246 -3480 253
rect -4473 219 -4466 225
rect -4484 208 -4477 215
rect -4284 209 -4278 216
rect -4225 209 -4219 216
rect -3112 425 -3106 433
rect -3026 429 -3020 436
rect -2945 422 -2936 430
rect -3031 340 -3023 349
rect -2967 340 -2961 348
rect -3103 322 -3098 329
rect -2966 249 -2960 256
rect -4092 199 -4084 207
rect -4127 187 -4119 196
rect -4671 175 -4663 183
rect -4532 172 -4524 178
rect -3953 176 -3947 183
rect -3894 176 -3888 183
rect -3638 176 -3632 183
rect -3579 176 -3573 183
rect -4541 157 -4536 163
rect -4365 134 -4360 141
rect -4304 134 -4298 141
rect -4198 133 -4191 138
rect -4224 120 -4219 128
rect -4501 109 -4494 116
rect -4462 79 -4455 86
rect -4671 68 -4663 76
rect -4541 57 -4536 63
rect -4671 -32 -4663 -24
rect -4034 101 -4029 108
rect -3973 101 -3967 108
rect -4072 84 -4066 92
rect -3867 100 -3860 105
rect -3719 101 -3714 108
rect -3658 101 -3652 108
rect -3893 87 -3888 95
rect -3552 100 -3545 105
rect -3578 87 -3573 95
rect -4370 45 -4364 53
rect -4284 49 -4278 56
rect -4203 42 -4194 50
rect -4289 -40 -4281 -31
rect -4225 -40 -4219 -32
rect -4361 -58 -4356 -51
rect -4254 -103 -4247 -95
rect -4223 -103 -4216 -95
rect -4092 -103 -4084 -95
rect -4039 12 -4033 20
rect -3953 16 -3947 23
rect -3872 9 -3863 17
rect -3958 -73 -3950 -64
rect -3894 -73 -3888 -65
rect -4030 -91 -4025 -84
rect -4072 -143 -4066 -136
rect -4484 -157 -4477 -149
rect -4284 -167 -4278 -160
rect -4225 -167 -4219 -160
rect -4501 -199 -4494 -194
rect -3923 -136 -3916 -128
rect -3724 12 -3718 20
rect -3638 16 -3632 23
rect -3557 9 -3548 17
rect -3643 -73 -3635 -64
rect -3579 -73 -3573 -65
rect -3715 -91 -3710 -84
rect -3578 -164 -3572 -157
rect -3678 -214 -3673 -209
rect -4541 -242 -4536 -235
rect -4365 -242 -4360 -235
rect -4304 -242 -4298 -235
rect -4198 -243 -4191 -238
rect -4224 -256 -4219 -248
rect -4515 -297 -4507 -290
rect -4370 -331 -4364 -323
rect -4284 -327 -4278 -320
rect -4203 -334 -4194 -326
rect -4289 -416 -4281 -407
rect -4225 -416 -4219 -408
rect -4361 -434 -4356 -427
rect -4254 -479 -4247 -471
<< metal2 >>
rect -4536 1606 -4407 1612
rect -4716 1517 -4670 1525
rect -4716 1425 -4708 1517
rect -4540 1512 -4536 1606
rect -4716 1417 -4670 1425
rect -4716 1318 -4708 1417
rect -4540 1405 -4536 1506
rect -4431 1482 -4425 1522
rect -4431 1476 -3813 1482
rect -4716 1310 -4670 1318
rect -4716 1218 -4708 1310
rect -4540 1305 -4536 1399
rect -4716 1210 -4670 1218
rect -4716 1115 -4708 1210
rect -4540 1202 -4536 1299
rect -4716 1107 -4670 1115
rect -4716 1015 -4708 1107
rect -4540 1102 -4536 1196
rect -4716 1007 -4670 1015
rect -4716 908 -4708 1007
rect -4540 995 -4536 1096
rect -4530 1052 -4524 1250
rect -4532 1044 -4524 1052
rect -4716 900 -4670 908
rect -4716 808 -4708 900
rect -4540 895 -4536 989
rect -4716 800 -4670 808
rect -4716 693 -4708 800
rect -4540 780 -4536 889
rect -4716 685 -4671 693
rect -4716 593 -4708 685
rect -4540 680 -4536 774
rect -4716 585 -4671 593
rect -4716 486 -4708 585
rect -4540 573 -4536 674
rect -4716 478 -4671 486
rect -4716 386 -4708 478
rect -4540 473 -4536 567
rect -4530 555 -4524 1044
rect -4520 673 -4512 1044
rect -4508 747 -4500 1350
rect -4496 1093 -4488 1457
rect -4297 1457 -4284 1464
rect -4219 1457 -3997 1464
rect -3932 1457 -3904 1464
rect -4297 1389 -4290 1457
rect -4393 1382 -4365 1389
rect -4298 1382 -4290 1389
rect -4393 1197 -4387 1382
rect -4297 1304 -4290 1382
rect -4198 1456 -4003 1457
rect -4198 1386 -4191 1456
rect -4010 1389 -4003 1456
rect -4105 1382 -4078 1389
rect -4011 1382 -4003 1389
rect -4224 1316 -4219 1368
rect -4224 1309 -4207 1316
rect -4297 1297 -4284 1304
rect -4213 1298 -4207 1309
rect -4370 1217 -4364 1293
rect -4213 1290 -4203 1298
rect -4370 1208 -4289 1217
rect -4203 1216 -4194 1290
rect -4219 1208 -4194 1216
rect -4105 1197 -4100 1382
rect -4010 1304 -4003 1382
rect -3911 1386 -3904 1457
rect -3937 1316 -3932 1368
rect -3937 1309 -3920 1316
rect -4010 1297 -3997 1304
rect -3926 1298 -3920 1309
rect -4083 1217 -4077 1293
rect -3926 1290 -3916 1298
rect -4083 1208 -4002 1217
rect -3916 1216 -3907 1290
rect -3932 1208 -3907 1216
rect -4393 1190 -4361 1197
rect -4105 1190 -4074 1197
rect -4247 1145 -4135 1153
rect -3820 1147 -3813 1476
rect -3809 1478 -3802 1486
rect -3809 1471 -3149 1478
rect -3665 1458 -3652 1465
rect -3587 1458 -3337 1465
rect -3272 1458 -3244 1465
rect -3665 1390 -3658 1458
rect -3761 1383 -3733 1390
rect -3666 1383 -3658 1390
rect -3761 1198 -3755 1383
rect -3665 1305 -3658 1383
rect -3566 1457 -3343 1458
rect -3566 1387 -3559 1457
rect -3350 1390 -3343 1457
rect -3445 1383 -3418 1390
rect -3351 1383 -3343 1390
rect -3592 1317 -3587 1369
rect -3592 1310 -3575 1317
rect -3665 1298 -3652 1305
rect -3581 1299 -3575 1310
rect -3738 1218 -3732 1294
rect -3581 1291 -3571 1299
rect -3738 1209 -3657 1218
rect -3571 1217 -3562 1291
rect -3587 1209 -3562 1217
rect -3445 1198 -3440 1383
rect -3350 1305 -3343 1383
rect -3251 1387 -3244 1458
rect -3277 1317 -3272 1369
rect -3277 1310 -3260 1317
rect -3350 1298 -3337 1305
rect -3266 1299 -3260 1310
rect -3423 1218 -3417 1294
rect -3266 1291 -3256 1299
rect -3423 1209 -3342 1218
rect -3256 1217 -3247 1291
rect -3272 1209 -3247 1217
rect -3761 1191 -3729 1198
rect -3445 1191 -3414 1198
rect -4143 1098 -4135 1145
rect -3953 1137 -3937 1144
rect -3828 1141 -3813 1147
rect -3615 1146 -3503 1154
rect -3953 1098 -3949 1137
rect -4143 1093 -3949 1098
rect -3945 1111 -3810 1115
rect -3945 1084 -3942 1111
rect -4032 1080 -3942 1084
rect -4297 1041 -4284 1048
rect -4219 1041 -3997 1048
rect -3932 1041 -3904 1048
rect -4297 973 -4290 1041
rect -4393 966 -4365 973
rect -4298 966 -4290 973
rect -4716 378 -4671 386
rect -4716 283 -4708 378
rect -4540 370 -4536 467
rect -4716 275 -4671 283
rect -4716 183 -4708 275
rect -4540 270 -4536 364
rect -4716 175 -4671 183
rect -4716 76 -4708 175
rect -4540 163 -4536 264
rect -4532 178 -4524 517
rect -4716 68 -4671 76
rect -4716 -24 -4708 68
rect -4540 63 -4536 157
rect -4716 -32 -4671 -24
rect -4541 -235 -4536 57
rect -4515 -290 -4507 418
rect -4496 304 -4489 944
rect -4485 602 -4477 726
rect -4473 225 -4466 627
rect -4501 -194 -4494 109
rect -4484 -149 -4477 208
rect -4462 86 -4455 841
rect -4393 781 -4387 966
rect -4297 888 -4290 966
rect -4198 1040 -4003 1041
rect -4198 970 -4191 1040
rect -4010 973 -4003 1040
rect -4105 966 -4078 973
rect -4011 966 -4003 973
rect -4224 900 -4219 952
rect -4224 893 -4207 900
rect -4297 881 -4284 888
rect -4213 882 -4207 893
rect -4370 801 -4364 877
rect -4213 874 -4203 882
rect -4370 792 -4289 801
rect -4203 800 -4194 874
rect -4219 792 -4194 800
rect -4105 781 -4100 966
rect -4010 888 -4003 966
rect -3911 970 -3904 1041
rect -3817 1047 -3810 1111
rect -3511 1090 -3503 1146
rect -3155 1147 -3149 1471
rect -3295 1138 -3277 1145
rect -3295 1090 -3290 1138
rect -3511 1083 -3290 1090
rect -3286 1110 -2876 1116
rect -3286 1079 -3281 1110
rect -3372 1073 -3281 1079
rect -3937 900 -3932 952
rect -3937 893 -3920 900
rect -4010 881 -3997 888
rect -3926 882 -3920 893
rect -4083 801 -4077 877
rect -3926 874 -3916 882
rect -4083 792 -4002 801
rect -3916 800 -3907 874
rect -3932 792 -3907 800
rect -4393 774 -4361 781
rect -4105 774 -4074 781
rect -4247 729 -4135 737
rect -4143 682 -4135 729
rect -3817 730 -3811 1047
rect -3664 1041 -3651 1048
rect -3586 1041 -3369 1048
rect -3304 1041 -3276 1048
rect -3664 973 -3657 1041
rect -3760 966 -3732 973
rect -3665 966 -3657 973
rect -3947 721 -3937 728
rect -3803 729 -3796 905
rect -3760 781 -3754 966
rect -3664 888 -3657 966
rect -3565 1040 -3375 1041
rect -3565 970 -3558 1040
rect -3382 973 -3375 1040
rect -3477 966 -3450 973
rect -3383 966 -3375 973
rect -3591 900 -3586 952
rect -3591 893 -3574 900
rect -3664 881 -3651 888
rect -3580 882 -3574 893
rect -3737 801 -3731 877
rect -3580 874 -3570 882
rect -3737 792 -3656 801
rect -3570 800 -3561 874
rect -3586 792 -3561 800
rect -3477 781 -3472 966
rect -3382 888 -3375 966
rect -3283 970 -3276 1041
rect -3309 900 -3304 952
rect -3309 893 -3292 900
rect -3382 881 -3369 888
rect -3298 882 -3292 893
rect -3455 801 -3449 877
rect -3298 874 -3288 882
rect -3455 792 -3374 801
rect -3288 800 -3279 874
rect -3304 792 -3279 800
rect -3760 774 -3728 781
rect -3477 774 -3446 781
rect -3614 729 -3502 737
rect -3947 682 -3940 721
rect -4143 675 -3940 682
rect -3510 684 -3502 729
rect -3188 731 -3181 1063
rect -3055 1046 -3042 1053
rect -2977 1046 -2949 1053
rect -3055 978 -3048 1046
rect -3153 971 -3123 978
rect -3056 971 -3048 978
rect -3153 786 -3145 971
rect -3055 893 -3048 971
rect -2956 975 -2949 1046
rect -2982 905 -2977 957
rect -2982 898 -2965 905
rect -3055 886 -3042 893
rect -2971 887 -2965 898
rect -3128 806 -3122 882
rect -2971 879 -2961 887
rect -3128 797 -3047 806
rect -2961 805 -2952 879
rect -2977 797 -2952 805
rect -3153 779 -3119 786
rect -2884 741 -2876 1110
rect -3005 734 -2876 741
rect -3320 721 -3309 728
rect -3320 684 -3313 721
rect -3510 677 -3313 684
rect -4297 583 -4284 590
rect -4219 583 -4191 590
rect -4297 515 -4290 583
rect -4395 508 -4365 515
rect -4298 508 -4290 515
rect -4429 -149 -4421 319
rect -4395 323 -4387 508
rect -4297 430 -4290 508
rect -4198 512 -4191 583
rect -4224 442 -4219 494
rect -4224 435 -4207 442
rect -4297 423 -4284 430
rect -4213 424 -4207 435
rect -4370 343 -4364 419
rect -4213 416 -4203 424
rect -4370 334 -4289 343
rect -4203 342 -4194 416
rect -4219 334 -4194 342
rect -4395 316 -4361 323
rect -4126 279 -4118 663
rect -3691 602 -3686 657
rect -3998 583 -3985 590
rect -3920 583 -3670 590
rect -3605 583 -3577 590
rect -3998 515 -3991 583
rect -4094 508 -4066 515
rect -3999 508 -3991 515
rect -4094 323 -4088 508
rect -3998 430 -3991 508
rect -3899 582 -3676 583
rect -3899 512 -3892 582
rect -3683 515 -3676 582
rect -3778 508 -3751 515
rect -3684 508 -3676 515
rect -3925 442 -3920 494
rect -3925 435 -3908 442
rect -3998 423 -3985 430
rect -3914 424 -3908 435
rect -4071 343 -4065 419
rect -3914 416 -3904 424
rect -4071 334 -3990 343
rect -3904 342 -3895 416
rect -3920 334 -3895 342
rect -3778 323 -3773 508
rect -3683 430 -3676 508
rect -3584 512 -3577 583
rect -3610 442 -3605 494
rect -3610 435 -3593 442
rect -3683 423 -3670 430
rect -3599 424 -3593 435
rect -3756 343 -3750 419
rect -3599 416 -3589 424
rect -3756 334 -3675 343
rect -3589 342 -3580 416
rect -3605 334 -3580 342
rect -4094 316 -4062 323
rect -3778 316 -3747 323
rect -4247 271 -4223 279
rect -3948 271 -3836 279
rect -4297 209 -4284 216
rect -4219 209 -4191 216
rect -4297 141 -4290 209
rect -4395 134 -4365 141
rect -4298 134 -4290 141
rect -4395 -51 -4387 134
rect -4297 56 -4290 134
rect -4198 138 -4191 209
rect -3844 215 -3836 271
rect -3488 253 -3480 665
rect -3354 589 -3341 596
rect -3276 589 -3026 596
rect -2961 589 -2933 596
rect -3354 521 -3347 589
rect -3450 514 -3422 521
rect -3355 514 -3347 521
rect -3450 329 -3444 514
rect -3354 436 -3347 514
rect -3255 588 -3032 589
rect -3255 518 -3248 588
rect -3039 521 -3032 588
rect -3134 514 -3107 521
rect -3040 514 -3032 521
rect -3281 448 -3276 500
rect -3281 441 -3264 448
rect -3354 429 -3341 436
rect -3270 430 -3264 441
rect -3427 349 -3421 425
rect -3270 422 -3260 430
rect -3427 340 -3346 349
rect -3260 348 -3251 422
rect -3276 340 -3251 348
rect -3134 329 -3129 514
rect -3039 436 -3032 514
rect -2940 518 -2933 589
rect -2966 448 -2961 500
rect -2966 441 -2949 448
rect -3039 429 -3026 436
rect -2955 430 -2949 441
rect -3112 349 -3106 425
rect -2955 422 -2945 430
rect -3112 340 -3031 349
rect -2945 348 -2936 422
rect -2961 340 -2936 348
rect -3450 322 -3418 329
rect -3134 322 -3103 329
rect -3304 277 -3192 285
rect -3618 243 -3610 250
rect -3618 215 -3613 243
rect -3844 208 -3613 215
rect -3200 221 -3192 277
rect -2974 249 -2966 256
rect -2974 221 -2969 249
rect -3200 214 -2969 221
rect -4224 68 -4219 120
rect -4224 61 -4207 68
rect -4297 49 -4284 56
rect -4213 50 -4207 61
rect -4370 -31 -4364 45
rect -4213 42 -4203 50
rect -4370 -40 -4289 -31
rect -4203 -32 -4194 42
rect -4219 -40 -4194 -32
rect -4395 -58 -4361 -51
rect -4247 -103 -4223 -95
rect -4127 -149 -4119 187
rect -4092 -95 -4084 199
rect -3966 176 -3953 183
rect -3888 176 -3638 183
rect -3573 176 -3545 183
rect -3966 108 -3959 176
rect -4062 101 -4034 108
rect -3967 101 -3959 108
rect -4072 -136 -4066 84
rect -4062 -84 -4056 101
rect -3966 23 -3959 101
rect -3867 175 -3644 176
rect -3867 105 -3860 175
rect -3651 108 -3644 175
rect -3746 101 -3719 108
rect -3652 101 -3644 108
rect -3893 35 -3888 87
rect -3893 28 -3876 35
rect -3966 16 -3953 23
rect -3882 17 -3876 28
rect -4039 -64 -4033 12
rect -3882 9 -3872 17
rect -4039 -73 -3958 -64
rect -3872 -65 -3863 9
rect -3888 -73 -3863 -65
rect -3746 -84 -3741 101
rect -3651 23 -3644 101
rect -3552 105 -3545 176
rect -3578 35 -3573 87
rect -3578 28 -3561 35
rect -3651 16 -3638 23
rect -3567 17 -3561 28
rect -3724 -64 -3718 12
rect -3567 9 -3557 17
rect -3724 -73 -3643 -64
rect -3557 -65 -3548 9
rect -3573 -73 -3548 -65
rect -4062 -91 -4030 -84
rect -3746 -91 -3715 -84
rect -3916 -136 -3804 -128
rect -4429 -155 -4119 -149
rect -4297 -167 -4284 -160
rect -4219 -167 -4191 -160
rect -4297 -235 -4290 -167
rect -4395 -242 -4365 -235
rect -4298 -242 -4290 -235
rect -4395 -427 -4387 -242
rect -4297 -320 -4290 -242
rect -4198 -238 -4191 -167
rect -3812 -192 -3804 -136
rect -3586 -164 -3578 -157
rect -3586 -192 -3581 -164
rect -3812 -199 -3581 -192
rect -4224 -308 -4219 -256
rect -4224 -315 -4207 -308
rect -4297 -327 -4284 -320
rect -4213 -326 -4207 -315
rect -4370 -407 -4364 -331
rect -4213 -334 -4203 -326
rect -4370 -416 -4289 -407
rect -4203 -408 -4194 -334
rect -4219 -416 -4194 -408
rect -4395 -434 -4361 -427
rect -3678 -471 -3673 -214
rect -4247 -479 -3673 -471
use full_adder  full_adder_0
timestamp 1668811232
transform 1 0 -5095 0 1 1416
box 671 68 1308 442
<< labels >>
rlabel metal1 -4665 1606 -4544 1612 5 drain
rlabel metal1 -4670 1417 -4579 1425 1 Gnd
rlabel metal1 -4665 1506 -4544 1512 5 drain
rlabel metal1 -4670 1310 -4579 1318 1 Gnd
rlabel metal1 -4665 1399 -4544 1405 5 drain
rlabel metal1 -4665 1299 -4544 1305 5 drain
rlabel metal1 -4665 889 -4544 895 5 drain
rlabel metal1 -4670 800 -4579 808 1 Gnd
rlabel metal1 -4665 989 -4544 995 5 drain
rlabel metal1 -4670 900 -4579 908 1 Gnd
rlabel metal1 -4665 1096 -4544 1102 5 drain
rlabel metal1 -4670 1007 -4579 1015 1 Gnd
rlabel metal1 -4670 1107 -4579 1115 1 Gnd
rlabel metal1 -4671 275 -4580 283 1 Gnd
rlabel metal1 -4666 364 -4545 370 5 drain
rlabel metal1 -4671 175 -4580 183 1 Gnd
rlabel metal1 -4666 264 -4545 270 5 drain
rlabel metal1 -4671 68 -4580 76 1 Gnd
rlabel metal1 -4666 157 -4545 163 5 drain
rlabel metal1 -4671 -32 -4580 -24 1 Gnd
rlabel metal1 -4666 57 -4545 63 5 drain
rlabel metal1 -4666 467 -4545 473 5 drain
rlabel metal1 -4671 378 -4580 386 1 Gnd
rlabel metal1 -4666 567 -4545 573 5 drain
rlabel metal1 -4671 478 -4580 486 1 Gnd
rlabel metal1 -4666 674 -4545 680 5 drain
rlabel metal1 -4671 585 -4580 593 1 Gnd
rlabel metal1 -4666 774 -4545 780 5 drain
rlabel metal1 -4671 685 -4580 693 1 Gnd
rlabel metal1 -4670 1517 -4579 1525 1 Gnd
rlabel metal1 -4665 1196 -4544 1202 5 drain
rlabel metal1 -4670 1210 -4579 1218 1 Gnd
rlabel polysilicon -4628 1447 -4623 1455 1 A3
rlabel polysilicon -4628 1036 -4623 1044 1 A2
rlabel polysilicon -4629 614 -4624 622 1 A1
rlabel polysilicon -4629 204 -4624 212 1 A0
rlabel polysilicon -4656 1552 -4651 1560 1 B3
rlabel polysilicon -4656 1450 -4651 1458 1 B2
rlabel polysilicon -4656 1346 -4651 1354 1 B1
rlabel polysilicon -4656 1249 -4651 1257 1 B0
rlabel metal1 -4559 7 -4552 19 1 P0
rlabel metal1 -4365 508 -4300 515 5 drain
rlabel metal1 -4370 419 -4300 427 1 Gnd
rlabel metal1 -4203 416 -4133 424 1 Gnd
rlabel metal1 -4198 505 -4133 512 5 drain
rlabel metal1 -4365 134 -4300 141 5 drain
rlabel metal1 -4370 45 -4300 53 1 Gnd
rlabel metal1 -4203 42 -4133 50 1 Gnd
rlabel metal1 -4198 131 -4133 138 5 drain
rlabel metal1 -4365 1382 -4300 1389 5 drain
rlabel metal1 -4370 1293 -4300 1301 1 Gnd
rlabel metal1 -4203 1290 -4133 1298 1 Gnd
rlabel metal1 -4198 1379 -4133 1386 5 drain
rlabel metal1 -4078 1382 -4013 1389 5 drain
rlabel metal1 -4083 1293 -4013 1301 1 Gnd
rlabel metal1 -3916 1290 -3846 1298 1 Gnd
rlabel metal1 -3911 1379 -3846 1386 5 drain
rlabel metal1 -3566 1380 -3501 1387 5 drain
rlabel metal1 -3571 1291 -3501 1299 1 Gnd
rlabel metal1 -3738 1294 -3668 1302 1 Gnd
rlabel metal1 -3733 1383 -3668 1390 5 drain
rlabel metal1 -3251 1380 -3186 1387 5 drain
rlabel metal1 -3256 1291 -3186 1299 1 Gnd
rlabel metal1 -3423 1294 -3353 1302 1 Gnd
rlabel metal1 -3418 1383 -3353 1390 5 drain
rlabel metal1 -3202 1317 -3194 1341 1 P5
rlabel metal1 -3565 963 -3500 970 5 drain
rlabel metal1 -3570 874 -3500 882 1 Gnd
rlabel metal1 -3737 877 -3667 885 1 Gnd
rlabel metal1 -3450 966 -3385 973 5 drain
rlabel metal1 -3455 877 -3385 885 1 Gnd
rlabel metal1 -3288 874 -3218 882 1 Gnd
rlabel metal1 -3283 963 -3218 970 5 drain
rlabel metal1 -2907 905 -2899 929 1 P4
rlabel metal1 -3123 971 -3058 978 5 drain
rlabel metal1 -3128 882 -3058 890 1 Gnd
rlabel metal1 -2961 879 -2891 887 1 Gnd
rlabel metal1 -2956 968 -2891 975 5 drain
rlabel metal1 -4365 966 -4300 973 5 drain
rlabel metal1 -4370 877 -4300 885 1 Gnd
rlabel metal1 -4203 874 -4133 882 1 Gnd
rlabel metal1 -4198 963 -4133 970 5 drain
rlabel metal1 -4078 966 -4013 973 5 drain
rlabel metal1 -4083 877 -4013 885 1 Gnd
rlabel metal1 -3916 874 -3846 882 1 Gnd
rlabel metal1 -3911 963 -3846 970 5 drain
rlabel metal1 -3899 505 -3834 512 5 drain
rlabel metal1 -3904 416 -3834 424 1 Gnd
rlabel metal1 -4071 419 -4001 427 1 Gnd
rlabel metal1 -4066 508 -4001 515 5 drain
rlabel metal1 -3584 505 -3519 512 5 drain
rlabel metal1 -3589 416 -3519 424 1 Gnd
rlabel metal1 -3756 419 -3686 427 1 Gnd
rlabel metal1 -3751 508 -3686 515 5 drain
rlabel metal1 -4198 -245 -4133 -238 5 drain
rlabel metal1 -4203 -334 -4133 -326 1 Gnd
rlabel metal1 -4370 -331 -4300 -323 1 Gnd
rlabel metal1 -4365 -242 -4300 -235 5 drain
rlabel metal1 -3719 101 -3654 108 5 drain
rlabel metal1 -3724 12 -3654 20 1 Gnd
rlabel metal1 -3557 9 -3487 17 1 Gnd
rlabel metal1 -3552 98 -3487 105 5 drain
rlabel metal1 -4034 101 -3969 108 5 drain
rlabel metal1 -4039 12 -3969 20 1 Gnd
rlabel metal1 -3872 9 -3802 17 1 Gnd
rlabel metal1 -3867 98 -3802 105 5 drain
rlabel metal1 -4149 -308 -4141 -284 1 P1
rlabel metal1 -3107 514 -3042 521 5 drain
rlabel metal1 -3112 425 -3042 433 1 Gnd
rlabel metal1 -2945 422 -2875 430 1 Gnd
rlabel metal1 -2940 511 -2875 518 5 drain
rlabel metal1 -3422 514 -3357 521 5 drain
rlabel metal1 -3427 425 -3357 433 1 Gnd
rlabel metal1 -3260 422 -3190 430 1 Gnd
rlabel metal1 -3255 511 -3190 518 5 drain
rlabel metal1 -3503 35 -3495 59 1 P2
rlabel metal1 -3732 966 -3667 973 5 drain
rlabel metal1 -2891 448 -2883 472 1 P3
rlabel polysilicon -4037 1135 -4033 1141 1 f2
rlabel metal1 -3786 1233 -3784 1246 1 f5
rlabel metal1 -3690 1072 -3688 1085 1 f6
rlabel polysilicon -3376 1132 -3374 1145 1 f7
rlabel polysilicon -4022 804 -4022 822 1 f8
rlabel metal2 -3801 754 -3799 772 1 f9
rlabel polysilicon -3693 850 -3691 868 1 f10
rlabel metal1 -3138 889 -3136 907 1 f11
rlabel polysilicon -4105 461 -4098 463 1 f12
rlabel polysilicon -3697 355 -3694 359 1 f13
rlabel metal1 -3465 355 -3463 379 1 f14
rlabel metal1 -3380 189 -3378 213 1 f15
rlabel metal1 -3122 394 -3120 418 1 f16
rlabel polysilicon -3065 265 -3062 273 1 f17
rlabel metal1 -2847 300 -2844 308 7 f18
rlabel polysilicon -3677 -149 -3674 -141 1 f19
rlabel polysilicon -4355 1336 -4352 1351 1 A2B3
rlabel polysilicon -4310 1221 -4307 1236 1 A3B2
rlabel metal1 -4380 743 -4377 758 1 A3B1
rlabel polysilicon -4327 848 -4324 863 1 A2B2
rlabel polysilicon -4327 517 -4324 532 1 A3B0
rlabel polysilicon -4355 459 -4352 474 1 A2B1
rlabel polysilicon -4355 83 -4352 98 1 A2B0
rlabel polysilicon -4327 18 -4324 33 1 A1B1
rlabel polysilicon -3997 -20 -3994 -5 1 A0B2
rlabel polysilicon -4356 -292 -4353 -277 1 A1B0
rlabel polysilicon -4327 -360 -4324 -345 1 A0B1
rlabel polysilicon -4029 393 -4026 407 1 A1B2
rlabel space -3801 1724 -3793 1733 1 P6
rlabel space -3791 1533 -3787 1539 1 C5
<< end >>
