**
.include TSMC_180nm.txt

.option scale=0.09u
.global Gnd

*capacitor
Cout output gnd 1.5f

*sources
V1  drain gnd dc 1
VA  A gnd pulse 1 0 0 0.1n 0.1n 40n 80n
VB  B gnd pulse 0 1 0 0.1n 0.1n 80n 160n 

***
* pulse(V1 V2 TD TR TF PW PER
* V1 = the initial amplitude
* V2 = the pulse amplitude
* TD = the delay time in seconds
* TR = the rise time in seconds
* TF = the fall time in seconds
* PW = the pulse width in seconds
* PER = the period in seconds
***

M1000 output B b_w_n Gnd CMOSN w=9 l=5
+  ad=135 pd=48 as=207 ps=64
M1001 output A drain w_n37_1# CMOSP w=8 l=5
+  ad=184 pd=62 as=184 ps=78
M1002 b_w_n A Gnd Gnd CMOSN w=9 l=5
+  ad=0 pd=0 as=126 ps=46
M1003 drain B output w_n37_1# CMOSP w=8 l=5
+  ad=0 pd=0 as=0 ps=0
C0 w_n37_1# A 0.12fF
C1 w_n37_1# B 0.12fF
C2 w_n37_1# output 0.03fF
C3 B output 0.20fF
C4 w_n37_1# drain 0.08fF
.tran 0.01us 1us

*Control 
.control

run
plot v(A) v(output)+2 v(B)+4

***
meas tran delay_a_lh
+trig v(a) val =0.5 rise=1 targ v(output) val =0.5 fall =1
meas tran delay_a_hl
+trig v(a) val =0.5 fall=1 targ v(output) val =0.5 rise =1

meas tran delay_b_lh
+trig v(b) val =0.5 rise=1 targ v(output) val =0.5 fall =1
meas tran delay_b_hl
+trig v(b) val =0.5 fall=1 targ v(output) val =0.5 rise =1

echo delay_a_lh: "$&delay_a_lh" 
echo delay_a_hl: "$&delay_a_hl" 
echo delay_b_lh: "$&delay_b_lh" 
echo delay_b_hl: "$&delay_b_hl"

.endc

.end
