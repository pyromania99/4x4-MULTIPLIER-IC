magic
tech scmos
timestamp 1668035305
<< nwell >>
rect -19 77 49 97
rect -100 2 -32 22
rect 67 -1 135 19
rect -19 -83 49 -63
<< ntransistor >>
rect -4 34 1 43
rect 24 34 29 43
rect -85 -41 -80 -32
rect -57 -41 -52 -32
rect 82 -44 87 -35
rect 110 -44 115 -35
rect -4 -126 1 -117
rect 24 -126 29 -117
<< ptransistor >>
rect -4 83 1 91
rect 24 83 29 91
rect -85 8 -80 16
rect -57 8 -52 16
rect 82 5 87 13
rect 110 5 115 13
rect -4 -77 1 -69
rect 24 -77 29 -69
<< ndiffusion >>
rect -10 34 -4 43
rect 1 34 24 43
rect 29 34 36 43
rect -91 -41 -85 -32
rect -80 -41 -57 -32
rect -52 -41 -45 -32
rect 76 -44 82 -35
rect 87 -44 110 -35
rect 115 -44 122 -35
rect -10 -126 -4 -117
rect 1 -126 24 -117
rect 29 -126 36 -117
<< pdiffusion >>
rect -6 83 -4 91
rect 1 83 9 91
rect 16 83 24 91
rect 29 83 36 91
rect -87 8 -85 16
rect -80 8 -72 16
rect -65 8 -57 16
rect -52 8 -45 16
rect 80 5 82 13
rect 87 5 95 13
rect 102 5 110 13
rect 115 5 122 13
rect -6 -77 -4 -69
rect 1 -77 9 -69
rect 16 -77 24 -69
rect 29 -77 36 -69
<< ndcontact >>
rect 6 106 13 113
rect 27 106 34 113
rect -75 31 -68 38
rect -54 31 -47 38
rect -18 34 -10 43
rect 36 34 44 43
rect 92 28 99 35
rect 113 28 120 35
rect -99 -41 -91 -32
rect -45 -41 -37 -32
rect 6 -54 13 -47
rect 68 -44 76 -35
rect 122 -44 130 -35
rect 30 -54 37 -47
rect -18 -126 -10 -117
rect 36 -126 44 -117
<< pdcontact >>
rect -13 83 -6 91
rect 9 83 16 91
rect 36 83 43 91
rect -94 8 -87 16
rect -72 8 -65 16
rect -45 8 -38 16
rect 73 5 80 13
rect 95 5 102 13
rect 122 5 129 13
rect -13 -77 -6 -69
rect 9 -77 16 -69
rect 36 -77 43 -69
<< psubstratepcontact >>
rect -6 17 2 25
rect -87 -58 -79 -50
rect 80 -61 88 -53
rect -6 -143 2 -135
rect 22 -143 30 -135
<< polysilicon >>
rect -4 91 1 99
rect 24 91 29 99
rect -4 66 1 83
rect -85 61 -81 66
rect -10 61 1 66
rect -85 16 -80 61
rect -4 43 1 61
rect 24 43 29 83
rect 44 59 49 67
rect -4 31 1 34
rect -57 16 -52 24
rect -85 -32 -80 8
rect -57 -32 -52 8
rect 24 -8 29 34
rect 82 13 87 59
rect 110 13 115 21
rect -37 -16 29 -8
rect -85 -44 -80 -41
rect -57 -89 -52 -41
rect -4 -69 1 -61
rect 24 -69 29 -16
rect 82 -35 87 5
rect 110 -35 115 5
rect 130 -19 138 -11
rect 82 -47 87 -44
rect -57 -95 -53 -89
rect -4 -117 1 -77
rect 24 -117 29 -77
rect 110 -93 115 -44
rect 44 -101 115 -93
rect -4 -129 1 -126
rect 24 -129 29 -126
<< polycontact >>
rect -81 61 -77 66
rect -14 61 -10 66
rect 36 59 44 67
rect 49 59 56 67
rect 81 59 87 67
rect -45 -16 -37 -8
rect 122 -19 130 -11
rect -53 -95 -48 -89
rect -9 -95 -4 -89
rect 36 -101 44 -93
<< metal1 >>
rect -7 106 6 113
rect 13 106 27 113
rect 34 106 46 113
rect -13 91 -6 106
rect 36 91 43 106
rect 9 67 16 83
rect -77 61 -14 66
rect 9 59 36 67
rect 56 59 81 67
rect 36 43 44 59
rect -94 31 -75 38
rect -68 31 -54 38
rect -47 31 -33 38
rect -94 16 -87 31
rect -45 16 -38 31
rect -18 25 -10 34
rect 80 30 92 35
rect 73 28 92 30
rect 99 28 113 35
rect 120 28 138 35
rect -18 17 -6 25
rect 2 17 47 25
rect 73 13 80 28
rect 122 13 129 28
rect -72 -8 -65 8
rect -72 -16 -45 -8
rect -45 -32 -37 -16
rect 95 -11 102 5
rect 95 -19 122 -11
rect 122 -35 130 -19
rect -99 -50 -91 -41
rect -93 -58 -87 -50
rect -79 -58 -29 -50
rect -7 -54 6 -47
rect 13 -54 30 -47
rect 37 -54 52 -47
rect 68 -53 76 -44
rect -13 -69 -6 -54
rect 36 -69 43 -54
rect 77 -61 80 -53
rect 88 -61 138 -53
rect -48 -95 -9 -89
rect 9 -93 16 -77
rect 9 -101 36 -93
rect 36 -117 44 -101
rect -18 -134 -10 -126
rect -10 -143 -6 -135
rect 2 -143 22 -135
rect 30 -143 46 -135
<< m2contact >>
rect -13 106 -7 113
rect 46 106 52 113
rect -33 31 -27 38
rect 73 30 80 35
rect 47 17 52 25
rect -99 -58 -93 -50
rect -13 -54 -7 -47
rect 68 -61 77 -53
rect -18 -143 -10 -134
rect 46 -143 52 -135
<< metal2 >>
rect -26 106 -13 113
rect 52 106 80 113
rect -26 38 -19 106
rect -27 31 -19 38
rect -26 -47 -19 31
rect 73 35 80 106
rect 47 -35 52 17
rect 47 -42 64 -35
rect -26 -54 -13 -47
rect 58 -53 64 -42
rect -99 -134 -93 -58
rect 58 -61 68 -53
rect -99 -143 -18 -134
rect 68 -135 77 -61
rect 52 -143 77 -135
<< labels >>
rlabel metal1 -94 31 -29 38 5 drain
rlabel metal1 -99 -58 -29 -50 1 Gnd
rlabel polysilicon -85 -32 -80 2 1 A
rlabel polysilicon -57 -32 -52 2 1 B
rlabel metal1 68 -61 138 -53 1 Gnd
rlabel metal1 73 28 138 35 5 drain
rlabel metal1 122 -35 130 -11 1 output
<< end >>
