magic
tech scmos
timestamp 1668810242
<< nwell >>
rect 606 367 674 387
rect 525 292 593 312
rect 692 289 760 309
rect 606 207 674 227
rect 529 101 597 121
rect 614 101 659 121
<< ntransistor >>
rect 621 324 626 333
rect 649 324 654 333
rect 540 249 545 258
rect 568 249 573 258
rect 707 246 712 255
rect 735 246 740 255
rect 621 164 626 173
rect 649 164 654 173
rect 544 58 549 67
rect 572 58 577 67
rect 629 58 634 67
<< ptransistor >>
rect 621 373 626 381
rect 649 373 654 381
rect 540 298 545 306
rect 568 298 573 306
rect 707 295 712 303
rect 735 295 740 303
rect 621 213 626 221
rect 649 213 654 221
rect 544 107 549 115
rect 572 107 577 115
rect 629 107 634 115
<< ndiffusion >>
rect 615 324 621 333
rect 626 324 649 333
rect 654 324 661 333
rect 534 249 540 258
rect 545 249 568 258
rect 573 249 580 258
rect 701 246 707 255
rect 712 246 735 255
rect 740 246 747 255
rect 615 164 621 173
rect 626 164 649 173
rect 654 164 661 173
rect 538 58 544 67
rect 549 58 572 67
rect 577 58 584 67
rect 621 58 629 67
rect 634 58 642 67
<< pdiffusion >>
rect 619 373 621 381
rect 626 373 634 381
rect 641 373 649 381
rect 654 373 661 381
rect 538 298 540 306
rect 545 298 553 306
rect 560 298 568 306
rect 573 298 580 306
rect 705 295 707 303
rect 712 295 720 303
rect 727 295 735 303
rect 740 295 747 303
rect 619 213 621 221
rect 626 213 634 221
rect 641 213 649 221
rect 654 213 661 221
rect 542 107 544 115
rect 549 107 557 115
rect 564 107 572 115
rect 577 107 584 115
rect 627 107 629 115
rect 634 107 642 115
rect 649 107 651 115
<< ndcontact >>
rect 631 396 638 403
rect 652 396 659 403
rect 550 321 557 328
rect 571 321 578 328
rect 607 324 615 333
rect 661 324 669 333
rect 717 318 724 325
rect 738 318 745 325
rect 526 249 534 258
rect 580 249 588 258
rect 631 236 638 243
rect 693 246 701 255
rect 747 246 755 255
rect 655 236 662 243
rect 554 130 561 136
rect 575 130 582 136
rect 607 164 615 173
rect 661 164 669 173
rect 627 130 635 136
rect 645 130 654 136
rect 530 58 538 67
rect 584 58 592 67
rect 613 58 621 67
rect 642 58 649 67
<< pdcontact >>
rect 612 373 619 381
rect 634 373 641 381
rect 661 373 668 381
rect 531 298 538 306
rect 553 298 560 306
rect 580 298 587 306
rect 698 295 705 303
rect 720 295 727 303
rect 747 295 754 303
rect 612 213 619 221
rect 634 213 641 221
rect 661 213 668 221
rect 535 107 542 115
rect 557 107 564 115
rect 584 107 591 115
rect 620 107 627 115
rect 642 107 649 115
<< psubstratepcontact >>
rect 619 307 627 315
rect 538 232 546 240
rect 705 229 713 237
rect 619 147 627 155
rect 647 147 655 155
rect 542 41 550 49
rect 581 41 589 49
rect 621 41 630 49
rect 640 41 649 49
<< polysilicon >>
rect 621 381 626 389
rect 649 381 654 389
rect 621 356 626 373
rect 540 351 544 356
rect 615 351 626 356
rect 540 306 545 351
rect 621 333 626 351
rect 649 333 654 373
rect 669 349 674 357
rect 621 321 626 324
rect 568 306 573 314
rect 540 273 545 298
rect 521 266 545 273
rect 540 258 545 266
rect 568 258 573 298
rect 649 282 654 324
rect 707 303 712 349
rect 735 303 740 311
rect 588 274 654 282
rect 540 246 545 249
rect 568 201 573 249
rect 621 221 626 229
rect 649 221 654 274
rect 707 255 712 295
rect 735 255 740 295
rect 707 243 712 246
rect 568 184 572 201
rect 568 180 589 184
rect 585 128 589 180
rect 621 173 626 213
rect 649 173 654 213
rect 735 197 740 246
rect 669 189 740 197
rect 621 161 626 164
rect 649 161 654 164
rect 572 123 589 128
rect 544 115 549 123
rect 572 115 577 123
rect 629 115 634 123
rect 544 84 549 107
rect 521 77 549 84
rect 544 67 549 77
rect 572 67 577 107
rect 629 91 634 107
rect 592 83 634 91
rect 629 67 634 83
rect 544 55 549 58
rect 572 55 577 58
rect 629 54 634 58
<< polycontact >>
rect 544 351 548 356
rect 611 351 615 356
rect 661 349 669 357
rect 674 349 681 357
rect 706 349 712 357
rect 513 266 521 273
rect 580 274 588 282
rect 572 195 577 201
rect 616 195 621 201
rect 661 189 669 197
rect 513 77 521 84
rect 568 70 572 74
rect 584 83 592 91
<< metal1 >>
rect 618 396 631 403
rect 638 396 652 403
rect 659 396 671 403
rect 612 381 619 396
rect 661 381 668 396
rect 634 357 641 373
rect 548 351 611 356
rect 634 349 661 357
rect 681 349 706 357
rect 661 333 669 349
rect 536 321 550 328
rect 557 321 571 328
rect 578 321 592 328
rect 531 306 538 321
rect 580 306 587 321
rect 607 315 615 324
rect 705 320 717 325
rect 698 318 717 320
rect 724 318 738 325
rect 745 318 763 325
rect 607 307 619 315
rect 627 307 672 315
rect 698 303 705 318
rect 747 303 754 318
rect 553 282 560 298
rect 553 274 580 282
rect 513 100 521 266
rect 580 258 588 274
rect 720 279 727 295
rect 720 271 788 279
rect 747 270 788 271
rect 747 255 755 270
rect 526 240 534 249
rect 532 232 538 240
rect 546 232 596 240
rect 618 236 631 243
rect 638 236 655 243
rect 662 236 677 243
rect 693 237 701 246
rect 612 221 619 236
rect 661 221 668 236
rect 702 229 705 237
rect 713 229 788 237
rect 577 195 616 201
rect 634 197 641 213
rect 634 189 661 197
rect 661 173 669 189
rect 607 156 615 164
rect 615 147 619 155
rect 627 147 647 155
rect 655 147 671 155
rect 540 130 554 136
rect 561 130 575 136
rect 582 130 627 136
rect 635 130 645 136
rect 654 130 657 136
rect 540 129 542 130
rect 535 115 542 129
rect 584 115 591 130
rect 620 115 627 130
rect 472 93 521 100
rect 513 84 521 93
rect 557 91 564 107
rect 557 83 584 91
rect 472 70 568 74
rect 584 67 592 83
rect 642 67 649 107
rect 530 49 538 58
rect 613 49 621 58
rect 660 49 669 147
rect 538 41 542 49
rect 550 41 581 49
rect 589 41 621 49
rect 630 41 640 49
rect 649 41 660 49
<< m2contact >>
rect 612 396 618 403
rect 671 396 677 403
rect 531 321 536 328
rect 592 321 598 328
rect 698 320 705 325
rect 672 307 677 315
rect 526 232 532 240
rect 612 236 618 243
rect 693 229 702 237
rect 607 147 615 156
rect 671 147 677 155
rect 535 129 540 136
rect 530 41 538 49
rect 660 41 669 49
<< metal2 >>
rect 599 396 612 403
rect 677 396 705 403
rect 599 328 606 396
rect 501 321 531 328
rect 598 321 606 328
rect 501 136 509 321
rect 599 243 606 321
rect 698 325 705 396
rect 672 255 677 307
rect 672 248 689 255
rect 599 236 612 243
rect 683 237 689 248
rect 526 156 532 232
rect 683 229 693 237
rect 526 147 607 156
rect 693 155 702 229
rect 677 147 702 155
rect 501 129 535 136
<< labels >>
rlabel metal1 698 318 763 325 5 drain
rlabel metal1 693 229 763 237 1 Gnd
rlabel polysilicon 568 258 573 292 1 B
rlabel polysilicon 540 258 545 292 1 A
rlabel metal1 526 232 596 240 1 Gnd
rlabel metal1 531 321 596 328 5 drain
rlabel metal1 642 84 649 92 1 Carry
rlabel metal1 747 255 755 279 1 Sum
<< end >>
