**
.include TSMC_180nm.txt

.option scale=0.09u
.global Gnd

*capacitor
Cout output gnd 1.5f

*sources
V1  drain gnd dc 1
VA  A gnd pulse 1 0 0 0.1n 0.1n 40n 80n
VB  B gnd pulse 0 1 0 0.1n 0.1n 80n 160n 

***
* pulse(V1 V2 TD TR TF PW PER
* V1 = the initial amplitude
* V2 = the pulse amplitude
* TD = the delay time in seconds
* TR = the rise time in seconds
* TF = the fall time in seconds
* PW = the pulse width in seconds
* PER = the period in seconds
***

M1000 Gnd B a_n200_n35# Gnd CMOSN w=5 l=4
+  ad=175 pd=100 as=115 ps=56
M1001 a_n200_7# A drain w_n219_1# CMOSP w=9 l=4
+  ad=207 pd=64 as=162 ps=72
M1002 output a_n200_n35# drain w_n145_1# CMOSP w=9 l=5
+  ad=99 pd=40 as=0 ps=0
M1003 output a_n200_n35# Gnd Gnd CMOSN w=5 l=5
+  ad=55 pd=32 as=0 ps=0
M1004 a_n200_n35# B a_n200_7# w_n219_1# CMOSP w=9 l=4
+  ad=108 pd=42 as=0 ps=0
M1005 a_n200_n35# A Gnd Gnd CMOSN w=5 l=4
+  ad=0 pd=0 as=0 ps=0
C0 w_n219_1# a_n200_n35# 0.04fF
C1 w_n145_1# a_n200_n35# 0.11fF
C2 w_n145_1# output 0.04fF
C3 B a_n200_n35# 0.12fF
C4 w_n219_1# drain 0.04fF
C5 w_n219_1# A 0.09fF
C6 w_n145_1# drain 0.04fF
C7 w_n219_1# B 0.09fF
C8 Gnd Gnd 0.47fF
C9 a_n200_n35# Gnd 0.79fF
C10 B Gnd 0.29fF
C11 A Gnd 0.28fF
C12 drain Gnd 0.38fF
C13 w_n145_1# Gnd 0.53fF
C14 w_n219_1# Gnd 1.37fF

.tran 0.01us 1us

*Control 
.control

run
plot v(A) v(output)+2 v(B)+4

***
meas tran delay_a_lh
+trig v(a) val =0.5 rise=1 targ v(output) val =0.5 fall =1
meas tran delay_a_hl
+trig v(a) val =0.5 fall=1 targ v(output) val =0.5 rise =1

meas tran delay_b_lh
+trig v(b) val =0.5 rise=1 targ v(output) val =0.5 fall =1
meas tran delay_b_hl
+trig v(b) val =0.5 fall=1 targ v(output) val =0.5 rise =1

echo delay_a_lh: "$&delay_a_lh" 
echo delay_a_hl: "$&delay_a_hl" 
echo delay_b_lh: "$&delay_b_lh" 
echo delay_b_hl: "$&delay_b_hl"

.endc

.end
