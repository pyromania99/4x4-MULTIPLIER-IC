magic
tech scmos
timestamp 1668810005
<< nwell >>
rect 790 405 858 425
rect 1105 405 1173 425
rect 709 330 777 350
rect 876 327 944 347
rect 1024 330 1092 350
rect 1191 327 1259 347
rect 790 245 858 265
rect 1105 245 1173 265
rect 713 139 781 159
rect 798 139 843 159
rect 1028 139 1096 159
rect 1113 139 1158 159
rect 1175 133 1239 154
rect 1248 133 1287 154
<< ntransistor >>
rect 805 362 810 371
rect 833 362 838 371
rect 1120 362 1125 371
rect 1148 362 1153 371
rect 724 287 729 296
rect 752 287 757 296
rect 891 284 896 293
rect 919 284 924 293
rect 1039 287 1044 296
rect 1067 287 1072 296
rect 1206 284 1211 293
rect 1234 284 1239 293
rect 805 202 810 211
rect 833 202 838 211
rect 1120 202 1125 211
rect 1148 202 1153 211
rect 728 96 733 105
rect 756 96 761 105
rect 813 96 818 105
rect 1043 96 1048 105
rect 1071 96 1076 105
rect 1128 96 1133 105
rect 1189 97 1193 102
rect 1216 97 1220 102
rect 1264 97 1269 102
<< ptransistor >>
rect 805 411 810 419
rect 833 411 838 419
rect 1120 411 1125 419
rect 1148 411 1153 419
rect 724 336 729 344
rect 752 336 757 344
rect 891 333 896 341
rect 919 333 924 341
rect 1039 336 1044 344
rect 1067 336 1072 344
rect 1206 333 1211 341
rect 1234 333 1239 341
rect 805 251 810 259
rect 833 251 838 259
rect 1120 251 1125 259
rect 1148 251 1153 259
rect 728 145 733 153
rect 756 145 761 153
rect 813 145 818 153
rect 1043 145 1048 153
rect 1071 145 1076 153
rect 1128 145 1133 153
rect 1189 139 1193 148
rect 1216 139 1220 148
rect 1264 139 1269 148
<< ndiffusion >>
rect 799 362 805 371
rect 810 362 833 371
rect 838 362 845 371
rect 1114 362 1120 371
rect 1125 362 1148 371
rect 1153 362 1160 371
rect 718 287 724 296
rect 729 287 752 296
rect 757 287 764 296
rect 885 284 891 293
rect 896 284 919 293
rect 924 284 931 293
rect 1033 287 1039 296
rect 1044 287 1067 296
rect 1072 287 1079 296
rect 1200 284 1206 293
rect 1211 284 1234 293
rect 1239 284 1246 293
rect 799 202 805 211
rect 810 202 833 211
rect 838 202 845 211
rect 1114 202 1120 211
rect 1125 202 1148 211
rect 1153 202 1160 211
rect 722 96 728 105
rect 733 96 756 105
rect 761 96 768 105
rect 805 96 813 105
rect 818 96 826 105
rect 1037 96 1043 105
rect 1048 96 1071 105
rect 1076 96 1083 105
rect 1120 96 1128 105
rect 1133 96 1141 105
rect 1185 97 1189 102
rect 1193 97 1200 102
rect 1206 97 1216 102
rect 1220 97 1226 102
rect 1255 97 1264 102
rect 1269 97 1275 102
<< pdiffusion >>
rect 803 411 805 419
rect 810 411 818 419
rect 825 411 833 419
rect 838 411 845 419
rect 1118 411 1120 419
rect 1125 411 1133 419
rect 1140 411 1148 419
rect 1153 411 1160 419
rect 722 336 724 344
rect 729 336 737 344
rect 744 336 752 344
rect 757 336 764 344
rect 889 333 891 341
rect 896 333 904 341
rect 911 333 919 341
rect 924 333 931 341
rect 1037 336 1039 344
rect 1044 336 1052 344
rect 1059 336 1067 344
rect 1072 336 1079 344
rect 1204 333 1206 341
rect 1211 333 1219 341
rect 1226 333 1234 341
rect 1239 333 1246 341
rect 803 251 805 259
rect 810 251 818 259
rect 825 251 833 259
rect 838 251 845 259
rect 1118 251 1120 259
rect 1125 251 1133 259
rect 1140 251 1148 259
rect 1153 251 1160 259
rect 726 145 728 153
rect 733 145 741 153
rect 748 145 756 153
rect 761 145 768 153
rect 811 145 813 153
rect 818 145 826 153
rect 833 145 835 153
rect 1041 145 1043 153
rect 1048 145 1056 153
rect 1063 145 1071 153
rect 1076 145 1083 153
rect 1126 145 1128 153
rect 1133 145 1141 153
rect 1148 145 1150 153
rect 1186 139 1189 148
rect 1193 139 1216 148
rect 1220 139 1227 148
rect 1259 139 1264 148
rect 1269 139 1275 148
<< ndcontact >>
rect 815 434 822 441
rect 836 434 843 441
rect 1130 434 1137 441
rect 1151 434 1158 441
rect 734 359 741 366
rect 755 359 762 366
rect 791 362 799 371
rect 845 362 853 371
rect 901 356 908 363
rect 922 356 929 363
rect 1049 359 1056 366
rect 1070 359 1077 366
rect 1106 362 1114 371
rect 1160 362 1168 371
rect 710 287 718 296
rect 764 287 772 296
rect 815 274 822 281
rect 1216 356 1223 363
rect 1237 356 1244 363
rect 877 284 885 293
rect 931 284 939 293
rect 1025 287 1033 296
rect 1079 287 1087 296
rect 839 274 846 281
rect 738 168 745 174
rect 759 168 766 174
rect 1130 274 1137 281
rect 1192 284 1200 293
rect 1246 284 1254 293
rect 1154 274 1161 281
rect 791 202 799 211
rect 845 202 853 211
rect 811 168 819 174
rect 829 168 838 174
rect 1053 168 1060 174
rect 1074 168 1081 174
rect 1106 202 1114 211
rect 1160 202 1168 211
rect 1126 168 1134 174
rect 1144 168 1153 174
rect 1190 163 1196 169
rect 1216 163 1222 169
rect 1243 163 1249 169
rect 1262 163 1268 169
rect 714 96 722 105
rect 768 96 776 105
rect 797 96 805 105
rect 826 96 833 105
rect 1029 96 1037 105
rect 1083 96 1091 105
rect 1112 96 1120 105
rect 1141 96 1148 105
rect 1180 97 1185 102
rect 1200 97 1206 102
rect 1226 97 1231 102
rect 1249 97 1255 102
rect 1275 97 1280 102
<< pdcontact >>
rect 796 411 803 419
rect 818 411 825 419
rect 845 411 852 419
rect 1111 411 1118 419
rect 1133 411 1140 419
rect 1160 411 1167 419
rect 715 336 722 344
rect 737 336 744 344
rect 764 336 771 344
rect 882 333 889 341
rect 904 333 911 341
rect 931 333 938 341
rect 1030 336 1037 344
rect 1052 336 1059 344
rect 1079 336 1086 344
rect 1197 333 1204 341
rect 1219 333 1226 341
rect 1246 333 1253 341
rect 796 251 803 259
rect 818 251 825 259
rect 845 251 852 259
rect 1111 251 1118 259
rect 1133 251 1140 259
rect 1160 251 1167 259
rect 719 145 726 153
rect 741 145 748 153
rect 768 145 775 153
rect 804 145 811 153
rect 826 145 833 153
rect 1034 145 1041 153
rect 1056 145 1063 153
rect 1083 145 1090 153
rect 1119 145 1126 153
rect 1141 145 1148 153
rect 1181 139 1186 148
rect 1227 139 1232 148
rect 1254 139 1259 148
rect 1275 139 1280 148
rect 1186 79 1192 85
rect 1217 79 1223 85
rect 1239 79 1245 85
rect 1258 79 1264 85
<< psubstratepcontact >>
rect 803 345 811 353
rect 1118 345 1126 353
rect 722 270 730 278
rect 889 267 897 275
rect 1037 270 1045 278
rect 1204 267 1212 275
rect 803 185 811 193
rect 831 185 839 193
rect 1118 185 1126 193
rect 1146 185 1154 193
rect 726 79 734 87
rect 805 79 814 87
rect 824 79 833 87
rect 1041 79 1049 87
rect 1120 79 1129 87
rect 1139 79 1148 87
<< polysilicon >>
rect 805 419 810 427
rect 833 419 838 427
rect 1120 419 1125 427
rect 1148 419 1153 427
rect 805 394 810 411
rect 724 389 728 394
rect 799 389 810 394
rect 724 344 729 389
rect 805 371 810 389
rect 833 371 838 411
rect 853 387 858 395
rect 1120 394 1125 411
rect 805 359 810 362
rect 752 344 757 352
rect 724 311 729 336
rect 705 304 729 311
rect 724 296 729 304
rect 752 296 757 336
rect 833 320 838 362
rect 891 341 896 387
rect 1039 389 1043 394
rect 1114 389 1125 394
rect 919 341 924 349
rect 1039 344 1044 389
rect 1120 371 1125 389
rect 1148 371 1153 411
rect 1168 387 1173 395
rect 1120 359 1125 362
rect 1067 344 1072 352
rect 772 312 838 320
rect 724 284 729 287
rect 752 239 757 287
rect 805 259 810 267
rect 833 259 838 312
rect 891 293 896 333
rect 919 293 924 333
rect 939 311 1020 317
rect 1039 311 1044 336
rect 939 309 1012 311
rect 1020 304 1044 311
rect 1039 296 1044 304
rect 1067 296 1072 336
rect 1148 320 1153 362
rect 1206 341 1211 387
rect 1234 341 1239 349
rect 1087 312 1153 320
rect 1039 284 1044 287
rect 891 281 896 284
rect 752 222 756 239
rect 752 218 773 222
rect 769 166 773 218
rect 805 211 810 251
rect 833 211 838 251
rect 919 235 924 284
rect 853 227 924 235
rect 1067 239 1072 287
rect 1120 259 1125 267
rect 1148 259 1153 312
rect 1206 293 1211 333
rect 1234 293 1239 333
rect 1206 281 1211 284
rect 1067 222 1071 239
rect 1067 218 1088 222
rect 805 199 810 202
rect 833 199 838 202
rect 1084 166 1088 218
rect 1120 211 1125 251
rect 1148 211 1153 251
rect 1234 235 1239 284
rect 1168 227 1239 235
rect 1120 199 1125 202
rect 1148 199 1153 202
rect 1164 170 1213 177
rect 756 161 773 166
rect 1071 161 1088 166
rect 728 153 733 161
rect 756 153 761 161
rect 813 153 818 161
rect 1043 153 1048 161
rect 1071 153 1076 161
rect 1128 153 1133 161
rect 728 122 733 145
rect 705 115 733 122
rect 728 105 733 115
rect 756 105 761 145
rect 813 129 818 145
rect 776 121 818 129
rect 1043 122 1048 145
rect 813 105 818 121
rect 1020 115 1048 122
rect 1043 105 1048 115
rect 1071 105 1076 145
rect 1128 129 1133 145
rect 1164 130 1168 170
rect 1207 160 1213 170
rect 1207 155 1220 160
rect 1189 148 1193 151
rect 1216 148 1220 155
rect 1264 148 1269 151
rect 1091 121 1133 129
rect 1153 123 1168 130
rect 1189 121 1193 139
rect 1128 105 1133 121
rect 1190 114 1193 121
rect 1189 102 1193 114
rect 1216 102 1220 139
rect 1264 119 1269 139
rect 1237 114 1269 119
rect 1264 102 1269 114
rect 728 93 733 96
rect 756 93 761 96
rect 813 92 818 96
rect 1043 93 1048 96
rect 1071 93 1076 96
rect 1128 92 1133 96
rect 1189 94 1193 97
rect 1216 93 1220 97
rect 1264 93 1269 97
<< polycontact >>
rect 728 389 732 394
rect 795 389 799 394
rect 845 387 853 395
rect 858 387 865 395
rect 890 387 896 395
rect 697 304 705 311
rect 1043 389 1047 394
rect 1110 389 1114 394
rect 1160 387 1168 395
rect 1173 387 1180 395
rect 1205 387 1211 395
rect 764 312 772 320
rect 931 309 939 317
rect 1012 304 1020 311
rect 1079 312 1087 320
rect 756 233 761 239
rect 800 233 805 239
rect 845 227 853 235
rect 1071 233 1076 239
rect 1115 233 1120 239
rect 1160 227 1168 235
rect 697 115 705 122
rect 752 108 756 112
rect 768 121 776 129
rect 1012 115 1020 122
rect 1083 121 1091 129
rect 1148 123 1153 130
rect 1183 114 1190 121
rect 1232 114 1237 119
<< metal1 >>
rect 802 434 815 441
rect 822 434 836 441
rect 843 434 855 441
rect 1117 434 1130 441
rect 1137 434 1151 441
rect 1158 434 1170 441
rect 796 419 803 434
rect 845 419 852 434
rect 1111 419 1118 434
rect 1160 419 1167 434
rect 818 395 825 411
rect 1133 395 1140 411
rect 732 389 795 394
rect 818 387 845 395
rect 865 387 890 395
rect 1047 389 1110 394
rect 1133 387 1160 395
rect 1180 387 1205 395
rect 845 371 853 387
rect 1160 371 1168 387
rect 720 359 734 366
rect 741 359 755 366
rect 762 359 776 366
rect 715 344 722 359
rect 764 344 771 359
rect 791 353 799 362
rect 889 358 901 363
rect 882 356 901 358
rect 908 356 922 363
rect 929 356 947 363
rect 1035 359 1049 366
rect 1056 359 1070 366
rect 1077 359 1091 366
rect 791 345 803 353
rect 811 345 856 353
rect 882 341 889 356
rect 931 341 938 356
rect 737 320 744 336
rect 1030 344 1037 359
rect 1079 344 1086 359
rect 1106 353 1114 362
rect 1204 358 1216 363
rect 1197 356 1216 358
rect 1223 356 1237 363
rect 1244 356 1274 363
rect 1106 345 1118 353
rect 1126 345 1171 353
rect 1197 341 1204 356
rect 1246 341 1253 356
rect 737 312 764 320
rect 697 205 705 304
rect 764 296 772 312
rect 904 317 911 333
rect 1052 320 1059 336
rect 904 309 931 317
rect 1052 312 1079 320
rect 931 293 939 309
rect 710 278 718 287
rect 716 270 722 278
rect 730 270 780 278
rect 802 274 815 281
rect 822 274 839 281
rect 846 274 861 281
rect 877 275 885 284
rect 796 259 803 274
rect 845 259 852 274
rect 886 267 889 275
rect 897 267 947 275
rect 761 233 800 239
rect 818 235 825 251
rect 818 227 845 235
rect 845 211 853 227
rect 671 200 705 205
rect 697 122 705 200
rect 791 194 799 202
rect 799 185 803 193
rect 811 185 831 193
rect 839 185 855 193
rect 724 168 738 174
rect 745 168 759 174
rect 766 168 811 174
rect 819 168 829 174
rect 838 168 841 174
rect 724 167 726 168
rect 719 153 726 167
rect 768 153 775 168
rect 804 153 811 168
rect 741 129 748 145
rect 741 121 768 129
rect 671 108 752 112
rect 768 105 776 121
rect 826 117 833 145
rect 826 105 833 109
rect 714 87 722 96
rect 797 87 805 96
rect 844 88 853 185
rect 1012 122 1020 304
rect 1079 296 1087 312
rect 1219 317 1226 333
rect 1219 309 1246 317
rect 1246 293 1254 308
rect 1025 278 1033 287
rect 1031 270 1037 278
rect 1045 270 1095 278
rect 1117 274 1130 281
rect 1137 274 1154 281
rect 1161 274 1176 281
rect 1192 275 1200 284
rect 1111 259 1118 274
rect 1160 259 1167 274
rect 1201 267 1204 275
rect 1212 267 1262 275
rect 1076 233 1115 239
rect 1133 235 1140 251
rect 1133 227 1160 235
rect 1160 211 1168 227
rect 1106 194 1114 202
rect 1114 185 1118 193
rect 1126 185 1146 193
rect 1154 185 1170 193
rect 1039 168 1053 174
rect 1060 168 1074 174
rect 1081 168 1126 174
rect 1134 168 1144 174
rect 1153 168 1156 174
rect 1039 167 1041 168
rect 1034 153 1041 167
rect 1083 153 1090 168
rect 1119 153 1126 168
rect 1056 129 1063 145
rect 1056 121 1083 129
rect 1083 105 1091 121
rect 1141 105 1148 145
rect 1029 88 1037 96
rect 844 87 1037 88
rect 1112 87 1120 96
rect 1159 87 1168 185
rect 1269 169 1274 356
rect 1181 163 1190 169
rect 1196 163 1216 169
rect 1222 163 1243 169
rect 1249 163 1262 169
rect 1268 163 1274 169
rect 1181 148 1186 163
rect 1254 148 1259 163
rect 1177 114 1183 121
rect 1227 119 1232 139
rect 1275 123 1280 139
rect 1200 114 1232 119
rect 1275 117 1308 123
rect 1200 102 1206 114
rect 1275 102 1280 117
rect 722 79 726 87
rect 734 79 805 87
rect 814 79 824 87
rect 833 79 1041 87
rect 1049 79 1120 87
rect 1129 79 1139 87
rect 1148 85 1168 87
rect 1180 85 1185 97
rect 1226 85 1231 97
rect 1249 85 1255 97
rect 1148 79 1186 85
rect 1192 79 1217 85
rect 1223 79 1239 85
rect 1245 79 1258 85
rect 1264 79 1268 85
<< m2contact >>
rect 796 434 802 441
rect 855 434 861 441
rect 1111 434 1117 441
rect 1170 434 1176 441
rect 715 359 720 366
rect 776 359 782 366
rect 882 358 889 363
rect 1030 359 1035 366
rect 1091 359 1097 366
rect 856 345 861 353
rect 1197 358 1204 363
rect 1171 345 1176 353
rect 710 270 716 278
rect 796 274 802 281
rect 877 267 886 275
rect 791 185 799 194
rect 855 185 861 193
rect 719 167 724 174
rect 826 109 833 117
rect 1246 308 1254 317
rect 1025 270 1031 278
rect 1111 274 1117 281
rect 1192 267 1201 275
rect 1106 185 1114 194
rect 1170 185 1176 193
rect 1034 167 1039 174
rect 1294 308 1302 317
rect 1171 114 1177 121
rect 714 79 722 87
rect 1268 79 1273 85
<< metal2 >>
rect 965 441 995 442
rect 783 434 796 441
rect 861 434 1111 441
rect 1176 434 1204 441
rect 783 366 790 434
rect 686 359 715 366
rect 782 359 790 366
rect 686 174 693 359
rect 783 281 790 359
rect 882 433 1105 434
rect 882 363 889 433
rect 1098 366 1105 433
rect 1003 359 1030 366
rect 1097 359 1105 366
rect 856 293 861 345
rect 856 286 873 293
rect 783 274 796 281
rect 867 275 873 286
rect 710 194 716 270
rect 867 267 877 275
rect 710 185 791 194
rect 877 193 886 267
rect 861 185 886 193
rect 1003 174 1008 359
rect 1098 281 1105 359
rect 1197 363 1204 434
rect 1171 293 1176 345
rect 1254 308 1294 317
rect 1171 286 1188 293
rect 1098 274 1111 281
rect 1182 275 1188 286
rect 1025 194 1031 270
rect 1182 267 1192 275
rect 1025 185 1106 194
rect 1192 193 1201 267
rect 1176 185 1201 193
rect 686 167 719 174
rect 1003 167 1034 174
rect 1160 117 1171 121
rect 833 114 1171 117
rect 833 109 1166 114
<< labels >>
rlabel metal1 882 356 947 363 5 drain
rlabel metal1 877 267 947 275 1 Gnd
rlabel metal1 710 270 780 278 1 Gnd
rlabel metal1 715 359 780 366 5 drain
rlabel polysilicon 724 296 729 330 1 A
rlabel polysilicon 752 296 757 330 1 B
rlabel metal1 1197 356 1262 363 5 drain
rlabel metal1 1192 267 1262 275 1 Gnd
rlabel metal1 1025 270 1095 278 1 Gnd
rlabel metal1 1030 359 1095 366 5 drain
rlabel metal1 1246 293 1254 317 1 Sum
rlabel polysilicon 1067 296 1072 330 1 Cin
rlabel metal1 931 293 939 317 1 S0
rlabel metal1 1141 122 1148 130 1 C1
rlabel metal1 1275 117 1280 125 1 C
rlabel m2contact 826 109 833 117 1 C0
<< end >>
