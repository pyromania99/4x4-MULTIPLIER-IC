magic
tech scmos
timestamp 1668813661
<< nwell >>
rect 132 346 200 366
rect 419 346 487 366
rect 51 271 119 291
rect 218 268 286 288
rect 338 271 406 291
rect 505 268 573 288
rect 132 186 200 206
rect 419 186 487 206
rect -249 92 -181 112
rect -164 92 -119 112
rect 55 80 123 100
rect 140 80 185 100
rect 342 80 410 100
rect 427 80 472 100
rect 489 74 553 95
rect 562 74 601 95
rect -249 -8 -181 12
rect -164 -8 -119 12
rect 132 -57 200 -37
rect 419 -57 487 -37
rect 764 -56 832 -36
rect 1079 -56 1147 -36
rect -249 -115 -181 -95
rect -164 -115 -119 -95
rect 51 -132 119 -112
rect 218 -135 286 -115
rect 338 -132 406 -112
rect 505 -135 573 -115
rect 683 -131 751 -111
rect 850 -134 918 -114
rect 998 -131 1066 -111
rect 1165 -134 1233 -114
rect -249 -215 -181 -195
rect -164 -215 -119 -195
rect 132 -217 200 -197
rect 419 -217 487 -197
rect 764 -216 832 -196
rect 1079 -216 1147 -196
rect -249 -318 -181 -298
rect -164 -318 -119 -298
rect 55 -323 123 -303
rect 140 -323 185 -303
rect 342 -323 410 -303
rect 427 -323 472 -303
rect 489 -329 553 -308
rect 562 -329 601 -308
rect 687 -322 755 -302
rect 772 -322 817 -302
rect 1002 -322 1070 -302
rect 1087 -322 1132 -302
rect 1149 -328 1213 -307
rect 1222 -328 1261 -307
rect -249 -418 -181 -398
rect -164 -418 -119 -398
rect 132 -473 200 -453
rect 419 -473 487 -453
rect 765 -473 833 -453
rect 1047 -473 1115 -453
rect 1374 -468 1442 -448
rect -249 -525 -181 -505
rect -164 -525 -119 -505
rect 51 -548 119 -528
rect 218 -551 286 -531
rect 338 -548 406 -528
rect 505 -551 573 -531
rect 684 -548 752 -528
rect 851 -551 919 -531
rect 966 -548 1034 -528
rect 1133 -551 1201 -531
rect 1293 -543 1361 -523
rect 1460 -546 1528 -526
rect -249 -625 -181 -605
rect -164 -625 -119 -605
rect 132 -633 200 -613
rect 419 -633 487 -613
rect 765 -633 833 -613
rect 1047 -633 1115 -613
rect 1374 -628 1442 -608
rect -250 -740 -182 -720
rect -165 -740 -120 -720
rect 55 -739 123 -719
rect 140 -739 185 -719
rect 342 -739 410 -719
rect 427 -739 472 -719
rect 489 -745 553 -724
rect 562 -745 601 -724
rect 688 -739 756 -719
rect 773 -739 818 -719
rect 970 -739 1038 -719
rect 1055 -739 1100 -719
rect 1117 -745 1181 -724
rect 1190 -745 1229 -724
rect 1297 -734 1365 -714
rect 1382 -734 1427 -714
rect -250 -840 -182 -820
rect -165 -840 -120 -820
rect -250 -947 -182 -927
rect -165 -947 -120 -927
rect 132 -931 200 -911
rect 431 -931 499 -911
rect 746 -931 814 -911
rect 1075 -925 1143 -905
rect 1390 -925 1458 -905
rect 51 -1006 119 -986
rect 218 -1009 286 -989
rect 350 -1006 418 -986
rect 517 -1009 585 -989
rect 665 -1006 733 -986
rect 832 -1009 900 -989
rect 994 -1000 1062 -980
rect 1161 -1003 1229 -983
rect 1309 -1000 1377 -980
rect 1476 -1003 1544 -983
rect -250 -1047 -182 -1027
rect -165 -1047 -120 -1027
rect 132 -1091 200 -1071
rect 431 -1091 499 -1071
rect 746 -1091 814 -1071
rect 1075 -1085 1143 -1065
rect 1390 -1085 1458 -1065
rect -250 -1150 -182 -1130
rect -165 -1150 -120 -1130
rect 55 -1197 123 -1177
rect 140 -1197 185 -1177
rect 354 -1197 422 -1177
rect 439 -1197 484 -1177
rect 669 -1197 737 -1177
rect 754 -1197 799 -1177
rect 998 -1191 1066 -1171
rect 1083 -1191 1128 -1171
rect 1313 -1191 1381 -1171
rect 1398 -1191 1443 -1171
rect 816 -1223 880 -1202
rect 889 -1223 928 -1202
rect 1460 -1217 1524 -1196
rect 1533 -1217 1572 -1196
rect -250 -1250 -182 -1230
rect -165 -1250 -120 -1230
rect 132 -1305 200 -1285
rect -250 -1357 -182 -1337
rect -165 -1357 -120 -1337
rect 463 -1338 531 -1318
rect 778 -1338 846 -1318
rect 51 -1380 119 -1360
rect 218 -1383 286 -1363
rect 382 -1413 450 -1393
rect 549 -1416 617 -1396
rect 697 -1413 765 -1393
rect 864 -1416 932 -1396
rect -250 -1457 -182 -1437
rect -165 -1457 -120 -1437
rect 132 -1465 200 -1445
rect 463 -1498 531 -1478
rect 778 -1498 846 -1478
rect 55 -1571 123 -1551
rect 140 -1571 185 -1551
rect 386 -1604 454 -1584
rect 471 -1604 516 -1584
rect 701 -1604 769 -1584
rect 786 -1604 831 -1584
rect 848 -1630 912 -1609
rect 921 -1630 960 -1609
rect 132 -1681 200 -1661
rect 51 -1756 119 -1736
rect 218 -1759 286 -1739
rect 132 -1841 200 -1821
rect 55 -1947 123 -1927
rect 140 -1947 185 -1927
<< ntransistor >>
rect 147 303 152 312
rect 175 303 180 312
rect 434 303 439 312
rect 462 303 467 312
rect 66 228 71 237
rect 94 228 99 237
rect 233 225 238 234
rect 261 225 266 234
rect 353 228 358 237
rect 381 228 386 237
rect 520 225 525 234
rect 548 225 553 234
rect 147 143 152 152
rect 175 143 180 152
rect 434 143 439 152
rect 462 143 467 152
rect -234 49 -229 58
rect -206 49 -201 58
rect -149 49 -144 58
rect 70 37 75 46
rect 98 37 103 46
rect 155 37 160 46
rect 357 37 362 46
rect 385 37 390 46
rect 442 37 447 46
rect 503 38 507 43
rect 530 38 534 43
rect 578 38 583 43
rect -234 -51 -229 -42
rect -206 -51 -201 -42
rect -149 -51 -144 -42
rect 147 -100 152 -91
rect 175 -100 180 -91
rect -234 -158 -229 -149
rect -206 -158 -201 -149
rect -149 -158 -144 -149
rect 434 -100 439 -91
rect 462 -100 467 -91
rect 66 -175 71 -166
rect 94 -175 99 -166
rect 779 -99 784 -90
rect 807 -99 812 -90
rect 233 -178 238 -169
rect 261 -178 266 -169
rect 353 -175 358 -166
rect 381 -175 386 -166
rect -234 -258 -229 -249
rect -206 -258 -201 -249
rect -149 -258 -144 -249
rect 1094 -99 1099 -90
rect 1122 -99 1127 -90
rect 520 -178 525 -169
rect 548 -178 553 -169
rect 698 -174 703 -165
rect 726 -174 731 -165
rect 147 -260 152 -251
rect 175 -260 180 -251
rect 865 -177 870 -168
rect 893 -177 898 -168
rect 1013 -174 1018 -165
rect 1041 -174 1046 -165
rect 434 -260 439 -251
rect 462 -260 467 -251
rect -234 -361 -229 -352
rect -206 -361 -201 -352
rect -149 -361 -144 -352
rect 1180 -177 1185 -168
rect 1208 -177 1213 -168
rect 779 -259 784 -250
rect 807 -259 812 -250
rect 1094 -259 1099 -250
rect 1122 -259 1127 -250
rect 70 -366 75 -357
rect 98 -366 103 -357
rect 155 -366 160 -357
rect 357 -366 362 -357
rect 385 -366 390 -357
rect 442 -366 447 -357
rect 503 -365 507 -360
rect 530 -365 534 -360
rect 578 -365 583 -360
rect 702 -365 707 -356
rect 730 -365 735 -356
rect 787 -365 792 -356
rect 1017 -365 1022 -356
rect 1045 -365 1050 -356
rect 1102 -365 1107 -356
rect 1163 -364 1167 -359
rect 1190 -364 1194 -359
rect 1238 -364 1243 -359
rect -234 -461 -229 -452
rect -206 -461 -201 -452
rect -149 -461 -144 -452
rect 147 -516 152 -507
rect 175 -516 180 -507
rect -234 -568 -229 -559
rect -206 -568 -201 -559
rect -149 -568 -144 -559
rect 434 -516 439 -507
rect 462 -516 467 -507
rect 66 -591 71 -582
rect 94 -591 99 -582
rect 780 -516 785 -507
rect 808 -516 813 -507
rect 233 -594 238 -585
rect 261 -594 266 -585
rect 353 -591 358 -582
rect 381 -591 386 -582
rect -234 -668 -229 -659
rect -206 -668 -201 -659
rect -149 -668 -144 -659
rect 1062 -516 1067 -507
rect 1090 -516 1095 -507
rect 520 -594 525 -585
rect 548 -594 553 -585
rect 699 -591 704 -582
rect 727 -591 732 -582
rect 147 -676 152 -667
rect 175 -676 180 -667
rect 1389 -511 1394 -502
rect 1417 -511 1422 -502
rect 866 -594 871 -585
rect 894 -594 899 -585
rect 981 -591 986 -582
rect 1009 -591 1014 -582
rect 434 -676 439 -667
rect 462 -676 467 -667
rect 1148 -594 1153 -585
rect 1176 -594 1181 -585
rect 1308 -586 1313 -577
rect 1336 -586 1341 -577
rect 780 -676 785 -667
rect 808 -676 813 -667
rect 1475 -589 1480 -580
rect 1503 -589 1508 -580
rect 1062 -676 1067 -667
rect 1090 -676 1095 -667
rect 1389 -671 1394 -662
rect 1417 -671 1422 -662
rect -235 -783 -230 -774
rect -207 -783 -202 -774
rect -150 -783 -145 -774
rect 70 -782 75 -773
rect 98 -782 103 -773
rect 155 -782 160 -773
rect 357 -782 362 -773
rect 385 -782 390 -773
rect 442 -782 447 -773
rect 503 -781 507 -776
rect 530 -781 534 -776
rect 578 -781 583 -776
rect 703 -782 708 -773
rect 731 -782 736 -773
rect 788 -782 793 -773
rect 985 -782 990 -773
rect 1013 -782 1018 -773
rect 1070 -782 1075 -773
rect 1131 -781 1135 -776
rect 1158 -781 1162 -776
rect 1206 -781 1211 -776
rect 1312 -777 1317 -768
rect 1340 -777 1345 -768
rect 1397 -777 1402 -768
rect -235 -883 -230 -874
rect -207 -883 -202 -874
rect -150 -883 -145 -874
rect -235 -990 -230 -981
rect -207 -990 -202 -981
rect -150 -990 -145 -981
rect 147 -974 152 -965
rect 175 -974 180 -965
rect 446 -974 451 -965
rect 474 -974 479 -965
rect 66 -1049 71 -1040
rect 94 -1049 99 -1040
rect -235 -1090 -230 -1081
rect -207 -1090 -202 -1081
rect -150 -1090 -145 -1081
rect 761 -974 766 -965
rect 789 -974 794 -965
rect 233 -1052 238 -1043
rect 261 -1052 266 -1043
rect 365 -1049 370 -1040
rect 393 -1049 398 -1040
rect 1090 -968 1095 -959
rect 1118 -968 1123 -959
rect 532 -1052 537 -1043
rect 560 -1052 565 -1043
rect 680 -1049 685 -1040
rect 708 -1049 713 -1040
rect 147 -1134 152 -1125
rect 175 -1134 180 -1125
rect 1405 -968 1410 -959
rect 1433 -968 1438 -959
rect 1009 -1043 1014 -1034
rect 1037 -1043 1042 -1034
rect 847 -1052 852 -1043
rect 875 -1052 880 -1043
rect 446 -1134 451 -1125
rect 474 -1134 479 -1125
rect 1176 -1046 1181 -1037
rect 1204 -1046 1209 -1037
rect 1324 -1043 1329 -1034
rect 1352 -1043 1357 -1034
rect 761 -1134 766 -1125
rect 789 -1134 794 -1125
rect 1491 -1046 1496 -1037
rect 1519 -1046 1524 -1037
rect 1090 -1128 1095 -1119
rect 1118 -1128 1123 -1119
rect 1405 -1128 1410 -1119
rect 1433 -1128 1438 -1119
rect -235 -1193 -230 -1184
rect -207 -1193 -202 -1184
rect -150 -1193 -145 -1184
rect 70 -1240 75 -1231
rect 98 -1240 103 -1231
rect 155 -1240 160 -1231
rect 369 -1240 374 -1231
rect 397 -1240 402 -1231
rect 454 -1240 459 -1231
rect 684 -1240 689 -1231
rect 712 -1240 717 -1231
rect 769 -1240 774 -1231
rect 1013 -1234 1018 -1225
rect 1041 -1234 1046 -1225
rect 1098 -1234 1103 -1225
rect 1328 -1234 1333 -1225
rect 1356 -1234 1361 -1225
rect 1413 -1234 1418 -1225
rect 830 -1259 834 -1254
rect 857 -1259 861 -1254
rect 905 -1259 910 -1254
rect 1474 -1253 1478 -1248
rect 1501 -1253 1505 -1248
rect 1549 -1253 1554 -1248
rect -235 -1293 -230 -1284
rect -207 -1293 -202 -1284
rect -150 -1293 -145 -1284
rect 147 -1348 152 -1339
rect 175 -1348 180 -1339
rect -235 -1400 -230 -1391
rect -207 -1400 -202 -1391
rect -150 -1400 -145 -1391
rect 66 -1423 71 -1414
rect 94 -1423 99 -1414
rect 478 -1381 483 -1372
rect 506 -1381 511 -1372
rect 233 -1426 238 -1417
rect 261 -1426 266 -1417
rect -235 -1500 -230 -1491
rect -207 -1500 -202 -1491
rect -150 -1500 -145 -1491
rect 793 -1381 798 -1372
rect 821 -1381 826 -1372
rect 397 -1456 402 -1447
rect 425 -1456 430 -1447
rect 147 -1508 152 -1499
rect 175 -1508 180 -1499
rect 564 -1459 569 -1450
rect 592 -1459 597 -1450
rect 712 -1456 717 -1447
rect 740 -1456 745 -1447
rect 879 -1459 884 -1450
rect 907 -1459 912 -1450
rect 478 -1541 483 -1532
rect 506 -1541 511 -1532
rect 793 -1541 798 -1532
rect 821 -1541 826 -1532
rect 70 -1614 75 -1605
rect 98 -1614 103 -1605
rect 155 -1614 160 -1605
rect 401 -1647 406 -1638
rect 429 -1647 434 -1638
rect 486 -1647 491 -1638
rect 716 -1647 721 -1638
rect 744 -1647 749 -1638
rect 801 -1647 806 -1638
rect 862 -1666 866 -1661
rect 889 -1666 893 -1661
rect 937 -1666 942 -1661
rect 147 -1724 152 -1715
rect 175 -1724 180 -1715
rect 66 -1799 71 -1790
rect 94 -1799 99 -1790
rect 233 -1802 238 -1793
rect 261 -1802 266 -1793
rect 147 -1884 152 -1875
rect 175 -1884 180 -1875
rect 70 -1990 75 -1981
rect 98 -1990 103 -1981
rect 155 -1990 160 -1981
<< ptransistor >>
rect 147 352 152 360
rect 175 352 180 360
rect 434 352 439 360
rect 462 352 467 360
rect 66 277 71 285
rect 94 277 99 285
rect 233 274 238 282
rect 261 274 266 282
rect 353 277 358 285
rect 381 277 386 285
rect 520 274 525 282
rect 548 274 553 282
rect 147 192 152 200
rect 175 192 180 200
rect 434 192 439 200
rect 462 192 467 200
rect -234 98 -229 106
rect -206 98 -201 106
rect -149 98 -144 106
rect 70 86 75 94
rect 98 86 103 94
rect 155 86 160 94
rect 357 86 362 94
rect 385 86 390 94
rect 442 86 447 94
rect 503 80 507 89
rect 530 80 534 89
rect 578 80 583 89
rect -234 -2 -229 6
rect -206 -2 -201 6
rect -149 -2 -144 6
rect 147 -51 152 -43
rect 175 -51 180 -43
rect 434 -51 439 -43
rect 462 -51 467 -43
rect 779 -50 784 -42
rect 807 -50 812 -42
rect 1094 -50 1099 -42
rect 1122 -50 1127 -42
rect -234 -109 -229 -101
rect -206 -109 -201 -101
rect -149 -109 -144 -101
rect 66 -126 71 -118
rect 94 -126 99 -118
rect 233 -129 238 -121
rect 261 -129 266 -121
rect 353 -126 358 -118
rect 381 -126 386 -118
rect -234 -209 -229 -201
rect -206 -209 -201 -201
rect -149 -209 -144 -201
rect 520 -129 525 -121
rect 548 -129 553 -121
rect 698 -125 703 -117
rect 726 -125 731 -117
rect 147 -211 152 -203
rect 175 -211 180 -203
rect 865 -128 870 -120
rect 893 -128 898 -120
rect 1013 -125 1018 -117
rect 1041 -125 1046 -117
rect 434 -211 439 -203
rect 462 -211 467 -203
rect 1180 -128 1185 -120
rect 1208 -128 1213 -120
rect 779 -210 784 -202
rect 807 -210 812 -202
rect -234 -312 -229 -304
rect -206 -312 -201 -304
rect -149 -312 -144 -304
rect 70 -317 75 -309
rect 98 -317 103 -309
rect 155 -317 160 -309
rect 357 -317 362 -309
rect 385 -317 390 -309
rect 442 -317 447 -309
rect 1094 -210 1099 -202
rect 1122 -210 1127 -202
rect 503 -323 507 -314
rect 530 -323 534 -314
rect 578 -323 583 -314
rect 702 -316 707 -308
rect 730 -316 735 -308
rect 787 -316 792 -308
rect 1017 -316 1022 -308
rect 1045 -316 1050 -308
rect 1102 -316 1107 -308
rect 1163 -322 1167 -313
rect 1190 -322 1194 -313
rect 1238 -322 1243 -313
rect -234 -412 -229 -404
rect -206 -412 -201 -404
rect -149 -412 -144 -404
rect 147 -467 152 -459
rect 175 -467 180 -459
rect 434 -467 439 -459
rect 462 -467 467 -459
rect 780 -467 785 -459
rect 808 -467 813 -459
rect 1062 -467 1067 -459
rect 1090 -467 1095 -459
rect 1389 -462 1394 -454
rect 1417 -462 1422 -454
rect -234 -519 -229 -511
rect -206 -519 -201 -511
rect -149 -519 -144 -511
rect 66 -542 71 -534
rect 94 -542 99 -534
rect 233 -545 238 -537
rect 261 -545 266 -537
rect 353 -542 358 -534
rect 381 -542 386 -534
rect -234 -619 -229 -611
rect -206 -619 -201 -611
rect -149 -619 -144 -611
rect 520 -545 525 -537
rect 548 -545 553 -537
rect 699 -542 704 -534
rect 727 -542 732 -534
rect 147 -627 152 -619
rect 175 -627 180 -619
rect 866 -545 871 -537
rect 894 -545 899 -537
rect 981 -542 986 -534
rect 1009 -542 1014 -534
rect 434 -627 439 -619
rect 462 -627 467 -619
rect 1308 -537 1313 -529
rect 1336 -537 1341 -529
rect 1148 -545 1153 -537
rect 1176 -545 1181 -537
rect 780 -627 785 -619
rect 808 -627 813 -619
rect -235 -734 -230 -726
rect -207 -734 -202 -726
rect -150 -734 -145 -726
rect 70 -733 75 -725
rect 98 -733 103 -725
rect 155 -733 160 -725
rect 357 -733 362 -725
rect 385 -733 390 -725
rect 442 -733 447 -725
rect 1475 -540 1480 -532
rect 1503 -540 1508 -532
rect 1062 -627 1067 -619
rect 1090 -627 1095 -619
rect 1389 -622 1394 -614
rect 1417 -622 1422 -614
rect 503 -739 507 -730
rect 530 -739 534 -730
rect 578 -739 583 -730
rect 703 -733 708 -725
rect 731 -733 736 -725
rect 788 -733 793 -725
rect 985 -733 990 -725
rect 1013 -733 1018 -725
rect 1070 -733 1075 -725
rect 1312 -728 1317 -720
rect 1340 -728 1345 -720
rect 1397 -728 1402 -720
rect 1131 -739 1135 -730
rect 1158 -739 1162 -730
rect 1206 -739 1211 -730
rect -235 -834 -230 -826
rect -207 -834 -202 -826
rect -150 -834 -145 -826
rect 147 -925 152 -917
rect 175 -925 180 -917
rect 446 -925 451 -917
rect 474 -925 479 -917
rect 761 -925 766 -917
rect 789 -925 794 -917
rect 1090 -919 1095 -911
rect 1118 -919 1123 -911
rect 1405 -919 1410 -911
rect 1433 -919 1438 -911
rect -235 -941 -230 -933
rect -207 -941 -202 -933
rect -150 -941 -145 -933
rect 66 -1000 71 -992
rect 94 -1000 99 -992
rect -235 -1041 -230 -1033
rect -207 -1041 -202 -1033
rect -150 -1041 -145 -1033
rect 233 -1003 238 -995
rect 261 -1003 266 -995
rect 365 -1000 370 -992
rect 393 -1000 398 -992
rect 532 -1003 537 -995
rect 560 -1003 565 -995
rect 680 -1000 685 -992
rect 708 -1000 713 -992
rect 147 -1085 152 -1077
rect 175 -1085 180 -1077
rect -235 -1144 -230 -1136
rect -207 -1144 -202 -1136
rect -150 -1144 -145 -1136
rect 1009 -994 1014 -986
rect 1037 -994 1042 -986
rect 847 -1003 852 -995
rect 875 -1003 880 -995
rect 446 -1085 451 -1077
rect 474 -1085 479 -1077
rect 1176 -997 1181 -989
rect 1204 -997 1209 -989
rect 1324 -994 1329 -986
rect 1352 -994 1357 -986
rect 761 -1085 766 -1077
rect 789 -1085 794 -1077
rect 1491 -997 1496 -989
rect 1519 -997 1524 -989
rect 1090 -1079 1095 -1071
rect 1118 -1079 1123 -1071
rect 1405 -1079 1410 -1071
rect 1433 -1079 1438 -1071
rect 70 -1191 75 -1183
rect 98 -1191 103 -1183
rect 155 -1191 160 -1183
rect 369 -1191 374 -1183
rect 397 -1191 402 -1183
rect 454 -1191 459 -1183
rect 684 -1191 689 -1183
rect 712 -1191 717 -1183
rect 769 -1191 774 -1183
rect 1013 -1185 1018 -1177
rect 1041 -1185 1046 -1177
rect 1098 -1185 1103 -1177
rect 1328 -1185 1333 -1177
rect 1356 -1185 1361 -1177
rect 1413 -1185 1418 -1177
rect 830 -1217 834 -1208
rect 857 -1217 861 -1208
rect 905 -1217 910 -1208
rect -235 -1244 -230 -1236
rect -207 -1244 -202 -1236
rect -150 -1244 -145 -1236
rect 1474 -1211 1478 -1202
rect 1501 -1211 1505 -1202
rect 1549 -1211 1554 -1202
rect 147 -1299 152 -1291
rect 175 -1299 180 -1291
rect -235 -1351 -230 -1343
rect -207 -1351 -202 -1343
rect -150 -1351 -145 -1343
rect 66 -1374 71 -1366
rect 94 -1374 99 -1366
rect 478 -1332 483 -1324
rect 506 -1332 511 -1324
rect 793 -1332 798 -1324
rect 821 -1332 826 -1324
rect 233 -1377 238 -1369
rect 261 -1377 266 -1369
rect -235 -1451 -230 -1443
rect -207 -1451 -202 -1443
rect -150 -1451 -145 -1443
rect 397 -1407 402 -1399
rect 425 -1407 430 -1399
rect 147 -1459 152 -1451
rect 175 -1459 180 -1451
rect 564 -1410 569 -1402
rect 592 -1410 597 -1402
rect 712 -1407 717 -1399
rect 740 -1407 745 -1399
rect 879 -1410 884 -1402
rect 907 -1410 912 -1402
rect 478 -1492 483 -1484
rect 506 -1492 511 -1484
rect 70 -1565 75 -1557
rect 98 -1565 103 -1557
rect 155 -1565 160 -1557
rect 793 -1492 798 -1484
rect 821 -1492 826 -1484
rect 401 -1598 406 -1590
rect 429 -1598 434 -1590
rect 486 -1598 491 -1590
rect 716 -1598 721 -1590
rect 744 -1598 749 -1590
rect 801 -1598 806 -1590
rect 862 -1624 866 -1615
rect 889 -1624 893 -1615
rect 937 -1624 942 -1615
rect 147 -1675 152 -1667
rect 175 -1675 180 -1667
rect 66 -1750 71 -1742
rect 94 -1750 99 -1742
rect 233 -1753 238 -1745
rect 261 -1753 266 -1745
rect 147 -1835 152 -1827
rect 175 -1835 180 -1827
rect 70 -1941 75 -1933
rect 98 -1941 103 -1933
rect 155 -1941 160 -1933
<< ndiffusion >>
rect 141 303 147 312
rect 152 303 175 312
rect 180 303 187 312
rect 428 303 434 312
rect 439 303 462 312
rect 467 303 474 312
rect 60 228 66 237
rect 71 228 94 237
rect 99 228 106 237
rect 227 225 233 234
rect 238 225 261 234
rect 266 225 273 234
rect 347 228 353 237
rect 358 228 381 237
rect 386 228 393 237
rect 514 225 520 234
rect 525 225 548 234
rect 553 225 560 234
rect 141 143 147 152
rect 152 143 175 152
rect 180 143 187 152
rect 428 143 434 152
rect 439 143 462 152
rect 467 143 474 152
rect -240 49 -234 58
rect -229 49 -206 58
rect -201 49 -194 58
rect -157 49 -149 58
rect -144 49 -136 58
rect 64 37 70 46
rect 75 37 98 46
rect 103 37 110 46
rect 147 37 155 46
rect 160 37 168 46
rect 351 37 357 46
rect 362 37 385 46
rect 390 37 397 46
rect 434 37 442 46
rect 447 37 455 46
rect 499 38 503 43
rect 507 38 514 43
rect 520 38 530 43
rect 534 38 540 43
rect 569 38 578 43
rect 583 38 589 43
rect -240 -51 -234 -42
rect -229 -51 -206 -42
rect -201 -51 -194 -42
rect -157 -51 -149 -42
rect -144 -51 -136 -42
rect 141 -100 147 -91
rect 152 -100 175 -91
rect 180 -100 187 -91
rect -240 -158 -234 -149
rect -229 -158 -206 -149
rect -201 -158 -194 -149
rect -157 -158 -149 -149
rect -144 -158 -136 -149
rect 428 -100 434 -91
rect 439 -100 462 -91
rect 467 -100 474 -91
rect 60 -175 66 -166
rect 71 -175 94 -166
rect 99 -175 106 -166
rect 773 -99 779 -90
rect 784 -99 807 -90
rect 812 -99 819 -90
rect 227 -178 233 -169
rect 238 -178 261 -169
rect 266 -178 273 -169
rect 347 -175 353 -166
rect 358 -175 381 -166
rect 386 -175 393 -166
rect -240 -258 -234 -249
rect -229 -258 -206 -249
rect -201 -258 -194 -249
rect -157 -258 -149 -249
rect -144 -258 -136 -249
rect 1088 -99 1094 -90
rect 1099 -99 1122 -90
rect 1127 -99 1134 -90
rect 514 -178 520 -169
rect 525 -178 548 -169
rect 553 -178 560 -169
rect 692 -174 698 -165
rect 703 -174 726 -165
rect 731 -174 738 -165
rect 141 -260 147 -251
rect 152 -260 175 -251
rect 180 -260 187 -251
rect 859 -177 865 -168
rect 870 -177 893 -168
rect 898 -177 905 -168
rect 1007 -174 1013 -165
rect 1018 -174 1041 -165
rect 1046 -174 1053 -165
rect 428 -260 434 -251
rect 439 -260 462 -251
rect 467 -260 474 -251
rect -240 -361 -234 -352
rect -229 -361 -206 -352
rect -201 -361 -194 -352
rect -157 -361 -149 -352
rect -144 -361 -136 -352
rect 1174 -177 1180 -168
rect 1185 -177 1208 -168
rect 1213 -177 1220 -168
rect 773 -259 779 -250
rect 784 -259 807 -250
rect 812 -259 819 -250
rect 1088 -259 1094 -250
rect 1099 -259 1122 -250
rect 1127 -259 1134 -250
rect 64 -366 70 -357
rect 75 -366 98 -357
rect 103 -366 110 -357
rect 147 -366 155 -357
rect 160 -366 168 -357
rect 351 -366 357 -357
rect 362 -366 385 -357
rect 390 -366 397 -357
rect 434 -366 442 -357
rect 447 -366 455 -357
rect 499 -365 503 -360
rect 507 -365 514 -360
rect 520 -365 530 -360
rect 534 -365 540 -360
rect 569 -365 578 -360
rect 583 -365 589 -360
rect 696 -365 702 -356
rect 707 -365 730 -356
rect 735 -365 742 -356
rect 779 -365 787 -356
rect 792 -365 800 -356
rect 1011 -365 1017 -356
rect 1022 -365 1045 -356
rect 1050 -365 1057 -356
rect 1094 -365 1102 -356
rect 1107 -365 1115 -356
rect 1159 -364 1163 -359
rect 1167 -364 1174 -359
rect 1180 -364 1190 -359
rect 1194 -364 1200 -359
rect 1229 -364 1238 -359
rect 1243 -364 1249 -359
rect -240 -461 -234 -452
rect -229 -461 -206 -452
rect -201 -461 -194 -452
rect -157 -461 -149 -452
rect -144 -461 -136 -452
rect 141 -516 147 -507
rect 152 -516 175 -507
rect 180 -516 187 -507
rect -240 -568 -234 -559
rect -229 -568 -206 -559
rect -201 -568 -194 -559
rect -157 -568 -149 -559
rect -144 -568 -136 -559
rect 428 -516 434 -507
rect 439 -516 462 -507
rect 467 -516 474 -507
rect 60 -591 66 -582
rect 71 -591 94 -582
rect 99 -591 106 -582
rect 774 -516 780 -507
rect 785 -516 808 -507
rect 813 -516 820 -507
rect 227 -594 233 -585
rect 238 -594 261 -585
rect 266 -594 273 -585
rect 347 -591 353 -582
rect 358 -591 381 -582
rect 386 -591 393 -582
rect -240 -668 -234 -659
rect -229 -668 -206 -659
rect -201 -668 -194 -659
rect -157 -668 -149 -659
rect -144 -668 -136 -659
rect 1056 -516 1062 -507
rect 1067 -516 1090 -507
rect 1095 -516 1102 -507
rect 514 -594 520 -585
rect 525 -594 548 -585
rect 553 -594 560 -585
rect 693 -591 699 -582
rect 704 -591 727 -582
rect 732 -591 739 -582
rect 141 -676 147 -667
rect 152 -676 175 -667
rect 180 -676 187 -667
rect 1383 -511 1389 -502
rect 1394 -511 1417 -502
rect 1422 -511 1429 -502
rect 860 -594 866 -585
rect 871 -594 894 -585
rect 899 -594 906 -585
rect 975 -591 981 -582
rect 986 -591 1009 -582
rect 1014 -591 1021 -582
rect 428 -676 434 -667
rect 439 -676 462 -667
rect 467 -676 474 -667
rect 1142 -594 1148 -585
rect 1153 -594 1176 -585
rect 1181 -594 1188 -585
rect 1302 -586 1308 -577
rect 1313 -586 1336 -577
rect 1341 -586 1348 -577
rect 774 -676 780 -667
rect 785 -676 808 -667
rect 813 -676 820 -667
rect 1469 -589 1475 -580
rect 1480 -589 1503 -580
rect 1508 -589 1515 -580
rect 1056 -676 1062 -667
rect 1067 -676 1090 -667
rect 1095 -676 1102 -667
rect 1383 -671 1389 -662
rect 1394 -671 1417 -662
rect 1422 -671 1429 -662
rect -241 -783 -235 -774
rect -230 -783 -207 -774
rect -202 -783 -195 -774
rect -158 -783 -150 -774
rect -145 -783 -137 -774
rect 64 -782 70 -773
rect 75 -782 98 -773
rect 103 -782 110 -773
rect 147 -782 155 -773
rect 160 -782 168 -773
rect 351 -782 357 -773
rect 362 -782 385 -773
rect 390 -782 397 -773
rect 434 -782 442 -773
rect 447 -782 455 -773
rect 499 -781 503 -776
rect 507 -781 514 -776
rect 520 -781 530 -776
rect 534 -781 540 -776
rect 569 -781 578 -776
rect 583 -781 589 -776
rect 697 -782 703 -773
rect 708 -782 731 -773
rect 736 -782 743 -773
rect 780 -782 788 -773
rect 793 -782 801 -773
rect 979 -782 985 -773
rect 990 -782 1013 -773
rect 1018 -782 1025 -773
rect 1062 -782 1070 -773
rect 1075 -782 1083 -773
rect 1127 -781 1131 -776
rect 1135 -781 1142 -776
rect 1148 -781 1158 -776
rect 1162 -781 1168 -776
rect 1197 -781 1206 -776
rect 1211 -781 1217 -776
rect 1306 -777 1312 -768
rect 1317 -777 1340 -768
rect 1345 -777 1352 -768
rect 1389 -777 1397 -768
rect 1402 -777 1410 -768
rect -241 -883 -235 -874
rect -230 -883 -207 -874
rect -202 -883 -195 -874
rect -158 -883 -150 -874
rect -145 -883 -137 -874
rect -241 -990 -235 -981
rect -230 -990 -207 -981
rect -202 -990 -195 -981
rect -158 -990 -150 -981
rect -145 -990 -137 -981
rect 141 -974 147 -965
rect 152 -974 175 -965
rect 180 -974 187 -965
rect 440 -974 446 -965
rect 451 -974 474 -965
rect 479 -974 486 -965
rect 60 -1049 66 -1040
rect 71 -1049 94 -1040
rect 99 -1049 106 -1040
rect -241 -1090 -235 -1081
rect -230 -1090 -207 -1081
rect -202 -1090 -195 -1081
rect -158 -1090 -150 -1081
rect -145 -1090 -137 -1081
rect 755 -974 761 -965
rect 766 -974 789 -965
rect 794 -974 801 -965
rect 227 -1052 233 -1043
rect 238 -1052 261 -1043
rect 266 -1052 273 -1043
rect 359 -1049 365 -1040
rect 370 -1049 393 -1040
rect 398 -1049 405 -1040
rect 1084 -968 1090 -959
rect 1095 -968 1118 -959
rect 1123 -968 1130 -959
rect 526 -1052 532 -1043
rect 537 -1052 560 -1043
rect 565 -1052 572 -1043
rect 674 -1049 680 -1040
rect 685 -1049 708 -1040
rect 713 -1049 720 -1040
rect 141 -1134 147 -1125
rect 152 -1134 175 -1125
rect 180 -1134 187 -1125
rect 1399 -968 1405 -959
rect 1410 -968 1433 -959
rect 1438 -968 1445 -959
rect 1003 -1043 1009 -1034
rect 1014 -1043 1037 -1034
rect 1042 -1043 1049 -1034
rect 841 -1052 847 -1043
rect 852 -1052 875 -1043
rect 880 -1052 887 -1043
rect 440 -1134 446 -1125
rect 451 -1134 474 -1125
rect 479 -1134 486 -1125
rect 1170 -1046 1176 -1037
rect 1181 -1046 1204 -1037
rect 1209 -1046 1216 -1037
rect 1318 -1043 1324 -1034
rect 1329 -1043 1352 -1034
rect 1357 -1043 1364 -1034
rect 755 -1134 761 -1125
rect 766 -1134 789 -1125
rect 794 -1134 801 -1125
rect 1485 -1046 1491 -1037
rect 1496 -1046 1519 -1037
rect 1524 -1046 1531 -1037
rect 1084 -1128 1090 -1119
rect 1095 -1128 1118 -1119
rect 1123 -1128 1130 -1119
rect 1399 -1128 1405 -1119
rect 1410 -1128 1433 -1119
rect 1438 -1128 1445 -1119
rect -241 -1193 -235 -1184
rect -230 -1193 -207 -1184
rect -202 -1193 -195 -1184
rect -158 -1193 -150 -1184
rect -145 -1193 -137 -1184
rect 64 -1240 70 -1231
rect 75 -1240 98 -1231
rect 103 -1240 110 -1231
rect 147 -1240 155 -1231
rect 160 -1240 168 -1231
rect 363 -1240 369 -1231
rect 374 -1240 397 -1231
rect 402 -1240 409 -1231
rect 446 -1240 454 -1231
rect 459 -1240 467 -1231
rect 678 -1240 684 -1231
rect 689 -1240 712 -1231
rect 717 -1240 724 -1231
rect 761 -1240 769 -1231
rect 774 -1240 782 -1231
rect 1007 -1234 1013 -1225
rect 1018 -1234 1041 -1225
rect 1046 -1234 1053 -1225
rect 1090 -1234 1098 -1225
rect 1103 -1234 1111 -1225
rect 1322 -1234 1328 -1225
rect 1333 -1234 1356 -1225
rect 1361 -1234 1368 -1225
rect 1405 -1234 1413 -1225
rect 1418 -1234 1426 -1225
rect 826 -1259 830 -1254
rect 834 -1259 841 -1254
rect 847 -1259 857 -1254
rect 861 -1259 867 -1254
rect 896 -1259 905 -1254
rect 910 -1259 916 -1254
rect 1470 -1253 1474 -1248
rect 1478 -1253 1485 -1248
rect 1491 -1253 1501 -1248
rect 1505 -1253 1511 -1248
rect 1540 -1253 1549 -1248
rect 1554 -1253 1560 -1248
rect -241 -1293 -235 -1284
rect -230 -1293 -207 -1284
rect -202 -1293 -195 -1284
rect -158 -1293 -150 -1284
rect -145 -1293 -137 -1284
rect 141 -1348 147 -1339
rect 152 -1348 175 -1339
rect 180 -1348 187 -1339
rect -241 -1400 -235 -1391
rect -230 -1400 -207 -1391
rect -202 -1400 -195 -1391
rect -158 -1400 -150 -1391
rect -145 -1400 -137 -1391
rect 60 -1423 66 -1414
rect 71 -1423 94 -1414
rect 99 -1423 106 -1414
rect 472 -1381 478 -1372
rect 483 -1381 506 -1372
rect 511 -1381 518 -1372
rect 227 -1426 233 -1417
rect 238 -1426 261 -1417
rect 266 -1426 273 -1417
rect -241 -1500 -235 -1491
rect -230 -1500 -207 -1491
rect -202 -1500 -195 -1491
rect -158 -1500 -150 -1491
rect -145 -1500 -137 -1491
rect 787 -1381 793 -1372
rect 798 -1381 821 -1372
rect 826 -1381 833 -1372
rect 391 -1456 397 -1447
rect 402 -1456 425 -1447
rect 430 -1456 437 -1447
rect 141 -1508 147 -1499
rect 152 -1508 175 -1499
rect 180 -1508 187 -1499
rect 558 -1459 564 -1450
rect 569 -1459 592 -1450
rect 597 -1459 604 -1450
rect 706 -1456 712 -1447
rect 717 -1456 740 -1447
rect 745 -1456 752 -1447
rect 873 -1459 879 -1450
rect 884 -1459 907 -1450
rect 912 -1459 919 -1450
rect 472 -1541 478 -1532
rect 483 -1541 506 -1532
rect 511 -1541 518 -1532
rect 787 -1541 793 -1532
rect 798 -1541 821 -1532
rect 826 -1541 833 -1532
rect 64 -1614 70 -1605
rect 75 -1614 98 -1605
rect 103 -1614 110 -1605
rect 147 -1614 155 -1605
rect 160 -1614 168 -1605
rect 395 -1647 401 -1638
rect 406 -1647 429 -1638
rect 434 -1647 441 -1638
rect 478 -1647 486 -1638
rect 491 -1647 499 -1638
rect 710 -1647 716 -1638
rect 721 -1647 744 -1638
rect 749 -1647 756 -1638
rect 793 -1647 801 -1638
rect 806 -1647 814 -1638
rect 858 -1666 862 -1661
rect 866 -1666 873 -1661
rect 879 -1666 889 -1661
rect 893 -1666 899 -1661
rect 928 -1666 937 -1661
rect 942 -1666 948 -1661
rect 141 -1724 147 -1715
rect 152 -1724 175 -1715
rect 180 -1724 187 -1715
rect 60 -1799 66 -1790
rect 71 -1799 94 -1790
rect 99 -1799 106 -1790
rect 227 -1802 233 -1793
rect 238 -1802 261 -1793
rect 266 -1802 273 -1793
rect 141 -1884 147 -1875
rect 152 -1884 175 -1875
rect 180 -1884 187 -1875
rect 64 -1990 70 -1981
rect 75 -1990 98 -1981
rect 103 -1990 110 -1981
rect 147 -1990 155 -1981
rect 160 -1990 168 -1981
<< pdiffusion >>
rect 145 352 147 360
rect 152 352 160 360
rect 167 352 175 360
rect 180 352 187 360
rect 432 352 434 360
rect 439 352 447 360
rect 454 352 462 360
rect 467 352 474 360
rect 64 277 66 285
rect 71 277 79 285
rect 86 277 94 285
rect 99 277 106 285
rect 231 274 233 282
rect 238 274 246 282
rect 253 274 261 282
rect 266 274 273 282
rect 351 277 353 285
rect 358 277 366 285
rect 373 277 381 285
rect 386 277 393 285
rect 518 274 520 282
rect 525 274 533 282
rect 540 274 548 282
rect 553 274 560 282
rect 145 192 147 200
rect 152 192 160 200
rect 167 192 175 200
rect 180 192 187 200
rect 432 192 434 200
rect 439 192 447 200
rect 454 192 462 200
rect 467 192 474 200
rect -236 98 -234 106
rect -229 98 -221 106
rect -214 98 -206 106
rect -201 98 -194 106
rect -151 98 -149 106
rect -144 98 -136 106
rect -129 98 -127 106
rect 68 86 70 94
rect 75 86 83 94
rect 90 86 98 94
rect 103 86 110 94
rect 153 86 155 94
rect 160 86 168 94
rect 175 86 177 94
rect 355 86 357 94
rect 362 86 370 94
rect 377 86 385 94
rect 390 86 397 94
rect 440 86 442 94
rect 447 86 455 94
rect 462 86 464 94
rect 500 80 503 89
rect 507 80 530 89
rect 534 80 541 89
rect 573 80 578 89
rect 583 80 589 89
rect -236 -2 -234 6
rect -229 -2 -221 6
rect -214 -2 -206 6
rect -201 -2 -194 6
rect -151 -2 -149 6
rect -144 -2 -136 6
rect -129 -2 -127 6
rect 145 -51 147 -43
rect 152 -51 160 -43
rect 167 -51 175 -43
rect 180 -51 187 -43
rect 432 -51 434 -43
rect 439 -51 447 -43
rect 454 -51 462 -43
rect 467 -51 474 -43
rect 777 -50 779 -42
rect 784 -50 792 -42
rect 799 -50 807 -42
rect 812 -50 819 -42
rect 1092 -50 1094 -42
rect 1099 -50 1107 -42
rect 1114 -50 1122 -42
rect 1127 -50 1134 -42
rect -236 -109 -234 -101
rect -229 -109 -221 -101
rect -214 -109 -206 -101
rect -201 -109 -194 -101
rect -151 -109 -149 -101
rect -144 -109 -136 -101
rect -129 -109 -127 -101
rect 64 -126 66 -118
rect 71 -126 79 -118
rect 86 -126 94 -118
rect 99 -126 106 -118
rect 231 -129 233 -121
rect 238 -129 246 -121
rect 253 -129 261 -121
rect 266 -129 273 -121
rect 351 -126 353 -118
rect 358 -126 366 -118
rect 373 -126 381 -118
rect 386 -126 393 -118
rect -236 -209 -234 -201
rect -229 -209 -221 -201
rect -214 -209 -206 -201
rect -201 -209 -194 -201
rect -151 -209 -149 -201
rect -144 -209 -136 -201
rect -129 -209 -127 -201
rect 518 -129 520 -121
rect 525 -129 533 -121
rect 540 -129 548 -121
rect 553 -129 560 -121
rect 696 -125 698 -117
rect 703 -125 711 -117
rect 718 -125 726 -117
rect 731 -125 738 -117
rect 145 -211 147 -203
rect 152 -211 160 -203
rect 167 -211 175 -203
rect 180 -211 187 -203
rect 863 -128 865 -120
rect 870 -128 878 -120
rect 885 -128 893 -120
rect 898 -128 905 -120
rect 1011 -125 1013 -117
rect 1018 -125 1026 -117
rect 1033 -125 1041 -117
rect 1046 -125 1053 -117
rect 432 -211 434 -203
rect 439 -211 447 -203
rect 454 -211 462 -203
rect 467 -211 474 -203
rect 1178 -128 1180 -120
rect 1185 -128 1193 -120
rect 1200 -128 1208 -120
rect 1213 -128 1220 -120
rect 777 -210 779 -202
rect 784 -210 792 -202
rect 799 -210 807 -202
rect 812 -210 819 -202
rect -236 -312 -234 -304
rect -229 -312 -221 -304
rect -214 -312 -206 -304
rect -201 -312 -194 -304
rect -151 -312 -149 -304
rect -144 -312 -136 -304
rect -129 -312 -127 -304
rect 68 -317 70 -309
rect 75 -317 83 -309
rect 90 -317 98 -309
rect 103 -317 110 -309
rect 153 -317 155 -309
rect 160 -317 168 -309
rect 175 -317 177 -309
rect 355 -317 357 -309
rect 362 -317 370 -309
rect 377 -317 385 -309
rect 390 -317 397 -309
rect 440 -317 442 -309
rect 447 -317 455 -309
rect 462 -317 464 -309
rect 1092 -210 1094 -202
rect 1099 -210 1107 -202
rect 1114 -210 1122 -202
rect 1127 -210 1134 -202
rect 500 -323 503 -314
rect 507 -323 530 -314
rect 534 -323 541 -314
rect 573 -323 578 -314
rect 583 -323 589 -314
rect 700 -316 702 -308
rect 707 -316 715 -308
rect 722 -316 730 -308
rect 735 -316 742 -308
rect 785 -316 787 -308
rect 792 -316 800 -308
rect 807 -316 809 -308
rect 1015 -316 1017 -308
rect 1022 -316 1030 -308
rect 1037 -316 1045 -308
rect 1050 -316 1057 -308
rect 1100 -316 1102 -308
rect 1107 -316 1115 -308
rect 1122 -316 1124 -308
rect 1160 -322 1163 -313
rect 1167 -322 1190 -313
rect 1194 -322 1201 -313
rect 1233 -322 1238 -313
rect 1243 -322 1249 -313
rect -236 -412 -234 -404
rect -229 -412 -221 -404
rect -214 -412 -206 -404
rect -201 -412 -194 -404
rect -151 -412 -149 -404
rect -144 -412 -136 -404
rect -129 -412 -127 -404
rect 145 -467 147 -459
rect 152 -467 160 -459
rect 167 -467 175 -459
rect 180 -467 187 -459
rect 432 -467 434 -459
rect 439 -467 447 -459
rect 454 -467 462 -459
rect 467 -467 474 -459
rect 778 -467 780 -459
rect 785 -467 793 -459
rect 800 -467 808 -459
rect 813 -467 820 -459
rect 1060 -467 1062 -459
rect 1067 -467 1075 -459
rect 1082 -467 1090 -459
rect 1095 -467 1102 -459
rect 1387 -462 1389 -454
rect 1394 -462 1402 -454
rect 1409 -462 1417 -454
rect 1422 -462 1429 -454
rect -236 -519 -234 -511
rect -229 -519 -221 -511
rect -214 -519 -206 -511
rect -201 -519 -194 -511
rect -151 -519 -149 -511
rect -144 -519 -136 -511
rect -129 -519 -127 -511
rect 64 -542 66 -534
rect 71 -542 79 -534
rect 86 -542 94 -534
rect 99 -542 106 -534
rect 231 -545 233 -537
rect 238 -545 246 -537
rect 253 -545 261 -537
rect 266 -545 273 -537
rect 351 -542 353 -534
rect 358 -542 366 -534
rect 373 -542 381 -534
rect 386 -542 393 -534
rect -236 -619 -234 -611
rect -229 -619 -221 -611
rect -214 -619 -206 -611
rect -201 -619 -194 -611
rect -151 -619 -149 -611
rect -144 -619 -136 -611
rect -129 -619 -127 -611
rect 518 -545 520 -537
rect 525 -545 533 -537
rect 540 -545 548 -537
rect 553 -545 560 -537
rect 697 -542 699 -534
rect 704 -542 712 -534
rect 719 -542 727 -534
rect 732 -542 739 -534
rect 145 -627 147 -619
rect 152 -627 160 -619
rect 167 -627 175 -619
rect 180 -627 187 -619
rect 864 -545 866 -537
rect 871 -545 879 -537
rect 886 -545 894 -537
rect 899 -545 906 -537
rect 979 -542 981 -534
rect 986 -542 994 -534
rect 1001 -542 1009 -534
rect 1014 -542 1021 -534
rect 432 -627 434 -619
rect 439 -627 447 -619
rect 454 -627 462 -619
rect 467 -627 474 -619
rect 1306 -537 1308 -529
rect 1313 -537 1321 -529
rect 1328 -537 1336 -529
rect 1341 -537 1348 -529
rect 1146 -545 1148 -537
rect 1153 -545 1161 -537
rect 1168 -545 1176 -537
rect 1181 -545 1188 -537
rect 778 -627 780 -619
rect 785 -627 793 -619
rect 800 -627 808 -619
rect 813 -627 820 -619
rect -237 -734 -235 -726
rect -230 -734 -222 -726
rect -215 -734 -207 -726
rect -202 -734 -195 -726
rect -152 -734 -150 -726
rect -145 -734 -137 -726
rect -130 -734 -128 -726
rect 68 -733 70 -725
rect 75 -733 83 -725
rect 90 -733 98 -725
rect 103 -733 110 -725
rect 153 -733 155 -725
rect 160 -733 168 -725
rect 175 -733 177 -725
rect 355 -733 357 -725
rect 362 -733 370 -725
rect 377 -733 385 -725
rect 390 -733 397 -725
rect 440 -733 442 -725
rect 447 -733 455 -725
rect 462 -733 464 -725
rect 1473 -540 1475 -532
rect 1480 -540 1488 -532
rect 1495 -540 1503 -532
rect 1508 -540 1515 -532
rect 1060 -627 1062 -619
rect 1067 -627 1075 -619
rect 1082 -627 1090 -619
rect 1095 -627 1102 -619
rect 1387 -622 1389 -614
rect 1394 -622 1402 -614
rect 1409 -622 1417 -614
rect 1422 -622 1429 -614
rect 500 -739 503 -730
rect 507 -739 530 -730
rect 534 -739 541 -730
rect 573 -739 578 -730
rect 583 -739 589 -730
rect 701 -733 703 -725
rect 708 -733 716 -725
rect 723 -733 731 -725
rect 736 -733 743 -725
rect 786 -733 788 -725
rect 793 -733 801 -725
rect 808 -733 810 -725
rect 983 -733 985 -725
rect 990 -733 998 -725
rect 1005 -733 1013 -725
rect 1018 -733 1025 -725
rect 1068 -733 1070 -725
rect 1075 -733 1083 -725
rect 1090 -733 1092 -725
rect 1310 -728 1312 -720
rect 1317 -728 1325 -720
rect 1332 -728 1340 -720
rect 1345 -728 1352 -720
rect 1395 -728 1397 -720
rect 1402 -728 1410 -720
rect 1417 -728 1419 -720
rect 1128 -739 1131 -730
rect 1135 -739 1158 -730
rect 1162 -739 1169 -730
rect 1201 -739 1206 -730
rect 1211 -739 1217 -730
rect -237 -834 -235 -826
rect -230 -834 -222 -826
rect -215 -834 -207 -826
rect -202 -834 -195 -826
rect -152 -834 -150 -826
rect -145 -834 -137 -826
rect -130 -834 -128 -826
rect 145 -925 147 -917
rect 152 -925 160 -917
rect 167 -925 175 -917
rect 180 -925 187 -917
rect 444 -925 446 -917
rect 451 -925 459 -917
rect 466 -925 474 -917
rect 479 -925 486 -917
rect 759 -925 761 -917
rect 766 -925 774 -917
rect 781 -925 789 -917
rect 794 -925 801 -917
rect 1088 -919 1090 -911
rect 1095 -919 1103 -911
rect 1110 -919 1118 -911
rect 1123 -919 1130 -911
rect 1403 -919 1405 -911
rect 1410 -919 1418 -911
rect 1425 -919 1433 -911
rect 1438 -919 1445 -911
rect -237 -941 -235 -933
rect -230 -941 -222 -933
rect -215 -941 -207 -933
rect -202 -941 -195 -933
rect -152 -941 -150 -933
rect -145 -941 -137 -933
rect -130 -941 -128 -933
rect 64 -1000 66 -992
rect 71 -1000 79 -992
rect 86 -1000 94 -992
rect 99 -1000 106 -992
rect -237 -1041 -235 -1033
rect -230 -1041 -222 -1033
rect -215 -1041 -207 -1033
rect -202 -1041 -195 -1033
rect -152 -1041 -150 -1033
rect -145 -1041 -137 -1033
rect -130 -1041 -128 -1033
rect 231 -1003 233 -995
rect 238 -1003 246 -995
rect 253 -1003 261 -995
rect 266 -1003 273 -995
rect 363 -1000 365 -992
rect 370 -1000 378 -992
rect 385 -1000 393 -992
rect 398 -1000 405 -992
rect 530 -1003 532 -995
rect 537 -1003 545 -995
rect 552 -1003 560 -995
rect 565 -1003 572 -995
rect 678 -1000 680 -992
rect 685 -1000 693 -992
rect 700 -1000 708 -992
rect 713 -1000 720 -992
rect 145 -1085 147 -1077
rect 152 -1085 160 -1077
rect 167 -1085 175 -1077
rect 180 -1085 187 -1077
rect -237 -1144 -235 -1136
rect -230 -1144 -222 -1136
rect -215 -1144 -207 -1136
rect -202 -1144 -195 -1136
rect -152 -1144 -150 -1136
rect -145 -1144 -137 -1136
rect -130 -1144 -128 -1136
rect 1007 -994 1009 -986
rect 1014 -994 1022 -986
rect 1029 -994 1037 -986
rect 1042 -994 1049 -986
rect 845 -1003 847 -995
rect 852 -1003 860 -995
rect 867 -1003 875 -995
rect 880 -1003 887 -995
rect 444 -1085 446 -1077
rect 451 -1085 459 -1077
rect 466 -1085 474 -1077
rect 479 -1085 486 -1077
rect 1174 -997 1176 -989
rect 1181 -997 1189 -989
rect 1196 -997 1204 -989
rect 1209 -997 1216 -989
rect 1322 -994 1324 -986
rect 1329 -994 1337 -986
rect 1344 -994 1352 -986
rect 1357 -994 1364 -986
rect 759 -1085 761 -1077
rect 766 -1085 774 -1077
rect 781 -1085 789 -1077
rect 794 -1085 801 -1077
rect 1489 -997 1491 -989
rect 1496 -997 1504 -989
rect 1511 -997 1519 -989
rect 1524 -997 1531 -989
rect 1088 -1079 1090 -1071
rect 1095 -1079 1103 -1071
rect 1110 -1079 1118 -1071
rect 1123 -1079 1130 -1071
rect 1403 -1079 1405 -1071
rect 1410 -1079 1418 -1071
rect 1425 -1079 1433 -1071
rect 1438 -1079 1445 -1071
rect 68 -1191 70 -1183
rect 75 -1191 83 -1183
rect 90 -1191 98 -1183
rect 103 -1191 110 -1183
rect 153 -1191 155 -1183
rect 160 -1191 168 -1183
rect 175 -1191 177 -1183
rect 367 -1191 369 -1183
rect 374 -1191 382 -1183
rect 389 -1191 397 -1183
rect 402 -1191 409 -1183
rect 452 -1191 454 -1183
rect 459 -1191 467 -1183
rect 474 -1191 476 -1183
rect 682 -1191 684 -1183
rect 689 -1191 697 -1183
rect 704 -1191 712 -1183
rect 717 -1191 724 -1183
rect 767 -1191 769 -1183
rect 774 -1191 782 -1183
rect 789 -1191 791 -1183
rect 1011 -1185 1013 -1177
rect 1018 -1185 1026 -1177
rect 1033 -1185 1041 -1177
rect 1046 -1185 1053 -1177
rect 1096 -1185 1098 -1177
rect 1103 -1185 1111 -1177
rect 1118 -1185 1120 -1177
rect 1326 -1185 1328 -1177
rect 1333 -1185 1341 -1177
rect 1348 -1185 1356 -1177
rect 1361 -1185 1368 -1177
rect 1411 -1185 1413 -1177
rect 1418 -1185 1426 -1177
rect 1433 -1185 1435 -1177
rect 827 -1217 830 -1208
rect 834 -1217 857 -1208
rect 861 -1217 868 -1208
rect 900 -1217 905 -1208
rect 910 -1217 916 -1208
rect -237 -1244 -235 -1236
rect -230 -1244 -222 -1236
rect -215 -1244 -207 -1236
rect -202 -1244 -195 -1236
rect -152 -1244 -150 -1236
rect -145 -1244 -137 -1236
rect -130 -1244 -128 -1236
rect 1471 -1211 1474 -1202
rect 1478 -1211 1501 -1202
rect 1505 -1211 1512 -1202
rect 1544 -1211 1549 -1202
rect 1554 -1211 1560 -1202
rect 145 -1299 147 -1291
rect 152 -1299 160 -1291
rect 167 -1299 175 -1291
rect 180 -1299 187 -1291
rect -237 -1351 -235 -1343
rect -230 -1351 -222 -1343
rect -215 -1351 -207 -1343
rect -202 -1351 -195 -1343
rect -152 -1351 -150 -1343
rect -145 -1351 -137 -1343
rect -130 -1351 -128 -1343
rect 64 -1374 66 -1366
rect 71 -1374 79 -1366
rect 86 -1374 94 -1366
rect 99 -1374 106 -1366
rect 476 -1332 478 -1324
rect 483 -1332 491 -1324
rect 498 -1332 506 -1324
rect 511 -1332 518 -1324
rect 791 -1332 793 -1324
rect 798 -1332 806 -1324
rect 813 -1332 821 -1324
rect 826 -1332 833 -1324
rect 231 -1377 233 -1369
rect 238 -1377 246 -1369
rect 253 -1377 261 -1369
rect 266 -1377 273 -1369
rect -237 -1451 -235 -1443
rect -230 -1451 -222 -1443
rect -215 -1451 -207 -1443
rect -202 -1451 -195 -1443
rect -152 -1451 -150 -1443
rect -145 -1451 -137 -1443
rect -130 -1451 -128 -1443
rect 395 -1407 397 -1399
rect 402 -1407 410 -1399
rect 417 -1407 425 -1399
rect 430 -1407 437 -1399
rect 145 -1459 147 -1451
rect 152 -1459 160 -1451
rect 167 -1459 175 -1451
rect 180 -1459 187 -1451
rect 562 -1410 564 -1402
rect 569 -1410 577 -1402
rect 584 -1410 592 -1402
rect 597 -1410 604 -1402
rect 710 -1407 712 -1399
rect 717 -1407 725 -1399
rect 732 -1407 740 -1399
rect 745 -1407 752 -1399
rect 877 -1410 879 -1402
rect 884 -1410 892 -1402
rect 899 -1410 907 -1402
rect 912 -1410 919 -1402
rect 476 -1492 478 -1484
rect 483 -1492 491 -1484
rect 498 -1492 506 -1484
rect 511 -1492 518 -1484
rect 68 -1565 70 -1557
rect 75 -1565 83 -1557
rect 90 -1565 98 -1557
rect 103 -1565 110 -1557
rect 153 -1565 155 -1557
rect 160 -1565 168 -1557
rect 175 -1565 177 -1557
rect 791 -1492 793 -1484
rect 798 -1492 806 -1484
rect 813 -1492 821 -1484
rect 826 -1492 833 -1484
rect 399 -1598 401 -1590
rect 406 -1598 414 -1590
rect 421 -1598 429 -1590
rect 434 -1598 441 -1590
rect 484 -1598 486 -1590
rect 491 -1598 499 -1590
rect 506 -1598 508 -1590
rect 714 -1598 716 -1590
rect 721 -1598 729 -1590
rect 736 -1598 744 -1590
rect 749 -1598 756 -1590
rect 799 -1598 801 -1590
rect 806 -1598 814 -1590
rect 821 -1598 823 -1590
rect 859 -1624 862 -1615
rect 866 -1624 889 -1615
rect 893 -1624 900 -1615
rect 932 -1624 937 -1615
rect 942 -1624 948 -1615
rect 145 -1675 147 -1667
rect 152 -1675 160 -1667
rect 167 -1675 175 -1667
rect 180 -1675 187 -1667
rect 64 -1750 66 -1742
rect 71 -1750 79 -1742
rect 86 -1750 94 -1742
rect 99 -1750 106 -1742
rect 231 -1753 233 -1745
rect 238 -1753 246 -1745
rect 253 -1753 261 -1745
rect 266 -1753 273 -1745
rect 145 -1835 147 -1827
rect 152 -1835 160 -1827
rect 167 -1835 175 -1827
rect 180 -1835 187 -1827
rect 68 -1941 70 -1933
rect 75 -1941 83 -1933
rect 90 -1941 98 -1933
rect 103 -1941 110 -1933
rect 153 -1941 155 -1933
rect 160 -1941 168 -1933
rect 175 -1941 177 -1933
<< ndcontact >>
rect 157 375 164 382
rect 178 375 185 382
rect 444 375 451 382
rect 465 375 472 382
rect 76 300 83 307
rect 97 300 104 307
rect 133 303 141 312
rect 187 303 195 312
rect 243 297 250 304
rect 264 297 271 304
rect 363 300 370 307
rect 387 300 394 307
rect 420 303 428 312
rect 474 303 482 312
rect 52 228 60 237
rect 106 228 114 237
rect 157 215 164 222
rect 530 297 537 304
rect 551 297 558 304
rect 219 225 227 234
rect 273 225 281 234
rect 339 228 347 237
rect 393 228 401 237
rect 181 215 188 222
rect -224 121 -217 127
rect -200 121 -193 127
rect -151 121 -143 127
rect -133 121 -124 127
rect 80 109 87 115
rect 101 109 108 115
rect 444 215 451 222
rect 506 225 514 234
rect 560 225 568 234
rect 468 215 475 222
rect 133 143 141 152
rect 187 143 195 152
rect 153 109 161 115
rect 171 109 180 115
rect 367 109 374 115
rect 388 109 395 115
rect 420 143 428 152
rect 474 143 482 152
rect 440 109 448 115
rect 458 109 467 115
rect -248 49 -240 58
rect -194 49 -186 58
rect -165 49 -157 58
rect -136 49 -129 58
rect -224 21 -217 27
rect 504 104 510 110
rect 530 104 536 110
rect 557 104 563 110
rect 576 104 582 110
rect 56 37 64 46
rect 110 37 118 46
rect 139 37 147 46
rect 168 37 175 46
rect 343 37 351 46
rect 397 37 405 46
rect 426 37 434 46
rect 455 37 462 46
rect 494 38 499 43
rect 514 38 520 43
rect 540 38 545 43
rect 563 38 569 43
rect 589 38 594 43
rect -197 21 -189 27
rect -151 21 -143 27
rect -133 21 -124 27
rect 157 -28 164 -21
rect 178 -28 185 -21
rect 444 -28 451 -21
rect 465 -28 472 -21
rect 789 -27 796 -20
rect 810 -27 817 -20
rect 1104 -27 1111 -20
rect 1125 -27 1132 -20
rect -248 -51 -240 -42
rect -194 -51 -186 -42
rect -165 -51 -157 -42
rect -136 -51 -129 -42
rect -224 -86 -217 -80
rect -151 -86 -143 -80
rect -133 -86 -124 -80
rect 76 -103 83 -96
rect 97 -103 104 -96
rect 133 -100 141 -91
rect 187 -100 195 -91
rect -248 -158 -240 -149
rect -194 -158 -186 -149
rect -165 -158 -157 -149
rect -136 -158 -129 -149
rect -224 -186 -217 -180
rect 243 -106 250 -99
rect 264 -106 271 -99
rect 363 -103 370 -96
rect 384 -103 391 -96
rect 420 -100 428 -91
rect 474 -100 482 -91
rect 52 -175 60 -166
rect 106 -175 114 -166
rect -197 -186 -190 -180
rect -151 -186 -143 -180
rect -133 -186 -124 -180
rect 157 -188 164 -181
rect 530 -106 537 -99
rect 551 -106 558 -99
rect 708 -102 715 -95
rect 729 -102 736 -95
rect 765 -99 773 -90
rect 819 -99 827 -90
rect 219 -178 227 -169
rect 273 -178 281 -169
rect 339 -175 347 -166
rect 393 -175 401 -166
rect 181 -188 188 -181
rect -248 -258 -240 -249
rect -194 -258 -186 -249
rect -165 -258 -157 -249
rect -136 -258 -129 -249
rect -224 -289 -217 -283
rect -201 -289 -194 -283
rect -151 -289 -143 -283
rect -133 -289 -124 -283
rect 80 -294 87 -288
rect 101 -294 108 -288
rect 444 -188 451 -181
rect 875 -105 882 -98
rect 896 -105 903 -98
rect 1023 -102 1030 -95
rect 1044 -102 1051 -95
rect 1080 -99 1088 -90
rect 1134 -99 1142 -90
rect 506 -178 514 -169
rect 560 -178 568 -169
rect 684 -174 692 -165
rect 738 -174 746 -165
rect 468 -188 475 -181
rect 133 -260 141 -251
rect 187 -260 195 -251
rect 153 -294 161 -288
rect 171 -294 180 -288
rect 367 -294 374 -288
rect 388 -294 395 -288
rect 789 -187 796 -180
rect 1190 -105 1197 -98
rect 1211 -105 1218 -98
rect 851 -177 859 -168
rect 905 -177 913 -168
rect 999 -174 1007 -165
rect 1053 -174 1061 -165
rect 813 -187 820 -180
rect 420 -260 428 -251
rect 474 -260 482 -251
rect 440 -294 448 -288
rect 458 -294 467 -288
rect -248 -361 -240 -352
rect -194 -361 -186 -352
rect -165 -361 -157 -352
rect -136 -361 -129 -352
rect 504 -299 510 -293
rect 712 -293 719 -287
rect 733 -293 740 -287
rect 530 -299 536 -293
rect 557 -299 563 -293
rect 576 -299 582 -293
rect 1104 -187 1111 -180
rect 1166 -177 1174 -168
rect 1220 -177 1228 -168
rect 1128 -187 1135 -180
rect 765 -259 773 -250
rect 819 -259 827 -250
rect 785 -293 793 -287
rect 803 -293 812 -287
rect 1027 -293 1034 -287
rect 1048 -293 1055 -287
rect 1080 -259 1088 -250
rect 1134 -259 1142 -250
rect 1100 -293 1108 -287
rect 1118 -293 1127 -287
rect -224 -389 -217 -383
rect 56 -366 64 -357
rect 110 -366 118 -357
rect 139 -366 147 -357
rect 168 -366 175 -357
rect 343 -366 351 -357
rect 397 -366 405 -357
rect 426 -366 434 -357
rect 455 -366 462 -357
rect 1164 -298 1170 -292
rect 1190 -298 1196 -292
rect 1217 -298 1223 -292
rect 1236 -298 1242 -292
rect 494 -365 499 -360
rect 514 -365 520 -360
rect 540 -365 545 -360
rect 563 -365 569 -360
rect 589 -365 594 -360
rect 688 -365 696 -356
rect 742 -365 750 -356
rect 771 -365 779 -356
rect 800 -365 807 -356
rect 1003 -365 1011 -356
rect 1057 -365 1065 -356
rect 1086 -365 1094 -356
rect 1115 -365 1122 -356
rect 1154 -364 1159 -359
rect 1174 -364 1180 -359
rect 1200 -364 1205 -359
rect 1223 -364 1229 -359
rect 1249 -364 1254 -359
rect -197 -389 -190 -383
rect -151 -389 -143 -383
rect -133 -389 -124 -383
rect 157 -444 164 -437
rect 178 -444 185 -437
rect 444 -444 451 -437
rect 465 -444 472 -437
rect 790 -444 797 -437
rect 811 -444 818 -437
rect 1072 -444 1079 -437
rect 1093 -444 1100 -437
rect 1399 -439 1406 -432
rect 1420 -439 1427 -432
rect -248 -461 -240 -452
rect -194 -461 -186 -452
rect -165 -461 -157 -452
rect -136 -461 -129 -452
rect -224 -496 -217 -490
rect -198 -496 -190 -490
rect -151 -496 -143 -490
rect -133 -496 -124 -490
rect 76 -519 83 -512
rect 97 -519 104 -512
rect 133 -516 141 -507
rect 187 -516 195 -507
rect -248 -568 -240 -559
rect -194 -568 -186 -559
rect -165 -568 -157 -559
rect -136 -568 -129 -559
rect -224 -596 -217 -590
rect 243 -522 250 -515
rect 264 -522 271 -515
rect 363 -519 370 -512
rect 384 -519 391 -512
rect 420 -516 428 -507
rect 474 -516 482 -507
rect -198 -596 -190 -590
rect -151 -596 -143 -590
rect -133 -596 -124 -590
rect 52 -591 60 -582
rect 106 -591 114 -582
rect 157 -604 164 -597
rect 530 -522 537 -515
rect 551 -522 558 -515
rect 709 -519 716 -512
rect 730 -519 737 -512
rect 766 -516 774 -507
rect 820 -516 828 -507
rect 219 -594 227 -585
rect 273 -594 281 -585
rect 339 -591 347 -582
rect 393 -591 401 -582
rect 181 -604 188 -597
rect -248 -668 -240 -659
rect -194 -668 -186 -659
rect -165 -668 -157 -659
rect -136 -668 -129 -659
rect -225 -711 -218 -705
rect -201 -711 -194 -705
rect -152 -711 -144 -705
rect -134 -711 -125 -705
rect 80 -710 87 -704
rect 101 -710 108 -704
rect 444 -604 451 -597
rect 876 -522 883 -515
rect 897 -522 904 -515
rect 991 -519 998 -512
rect 1012 -519 1019 -512
rect 1048 -516 1056 -507
rect 1102 -516 1110 -507
rect 506 -594 514 -585
rect 560 -594 568 -585
rect 685 -591 693 -582
rect 739 -591 747 -582
rect 468 -604 475 -597
rect 133 -676 141 -667
rect 187 -676 195 -667
rect 153 -710 161 -704
rect 171 -710 180 -704
rect 367 -710 374 -704
rect 388 -710 395 -704
rect 790 -604 797 -597
rect 1158 -522 1165 -515
rect 1179 -522 1186 -515
rect 1318 -514 1325 -507
rect 1339 -514 1346 -507
rect 1375 -511 1383 -502
rect 1429 -511 1437 -502
rect 852 -594 860 -585
rect 906 -594 914 -585
rect 967 -591 975 -582
rect 1021 -591 1029 -582
rect 814 -604 821 -597
rect 420 -676 428 -667
rect 474 -676 482 -667
rect 440 -710 448 -704
rect 458 -710 467 -704
rect 504 -715 510 -709
rect 530 -715 536 -709
rect 557 -715 563 -709
rect 576 -715 582 -709
rect 713 -710 720 -704
rect 734 -710 741 -704
rect 1072 -604 1079 -597
rect 1485 -517 1492 -510
rect 1506 -517 1513 -510
rect 1134 -594 1142 -585
rect 1188 -594 1196 -585
rect 1294 -586 1302 -577
rect 1348 -586 1356 -577
rect 1096 -604 1103 -597
rect 766 -676 774 -667
rect 820 -676 828 -667
rect 786 -710 794 -704
rect 804 -710 813 -704
rect 995 -710 1002 -704
rect 1016 -710 1023 -704
rect 1399 -599 1406 -592
rect 1461 -589 1469 -580
rect 1515 -589 1523 -580
rect 1423 -599 1430 -592
rect 1048 -676 1056 -667
rect 1102 -676 1110 -667
rect 1068 -710 1076 -704
rect 1086 -710 1095 -704
rect 1322 -705 1329 -699
rect 1343 -705 1350 -699
rect 1375 -671 1383 -662
rect 1429 -671 1437 -662
rect 1395 -705 1403 -699
rect 1413 -705 1422 -699
rect -249 -783 -241 -774
rect -195 -783 -187 -774
rect -166 -783 -158 -774
rect -137 -783 -130 -774
rect 56 -782 64 -773
rect 110 -782 118 -773
rect 139 -782 147 -773
rect 168 -782 175 -773
rect 343 -782 351 -773
rect 397 -782 405 -773
rect 426 -782 434 -773
rect 455 -782 462 -773
rect 1132 -715 1138 -709
rect 1158 -715 1164 -709
rect 1185 -715 1191 -709
rect 1204 -715 1210 -709
rect 494 -781 499 -776
rect 514 -781 520 -776
rect 540 -781 545 -776
rect 563 -781 569 -776
rect 589 -781 594 -776
rect -225 -811 -218 -805
rect -200 -811 -192 -805
rect -152 -811 -144 -805
rect -134 -811 -125 -805
rect 689 -782 697 -773
rect 743 -782 751 -773
rect 772 -782 780 -773
rect 801 -782 808 -773
rect 971 -782 979 -773
rect 1025 -782 1033 -773
rect 1054 -782 1062 -773
rect 1083 -782 1090 -773
rect 1122 -781 1127 -776
rect 1142 -781 1148 -776
rect 1168 -781 1173 -776
rect 1191 -781 1197 -776
rect 1217 -781 1222 -776
rect 1298 -777 1306 -768
rect 1352 -777 1360 -768
rect 1381 -777 1389 -768
rect 1410 -777 1417 -768
rect -249 -883 -241 -874
rect -195 -883 -187 -874
rect -166 -883 -158 -874
rect -137 -883 -130 -874
rect -225 -918 -218 -912
rect 157 -902 164 -895
rect 178 -902 185 -895
rect 456 -902 463 -895
rect 477 -902 484 -895
rect 771 -902 778 -895
rect 792 -902 799 -895
rect 1100 -896 1107 -889
rect 1121 -896 1128 -889
rect 1415 -896 1422 -889
rect 1436 -896 1443 -889
rect -200 -918 -193 -912
rect -152 -918 -144 -912
rect -134 -918 -125 -912
rect -249 -990 -241 -981
rect -195 -990 -187 -981
rect -166 -990 -158 -981
rect -137 -990 -130 -981
rect -225 -1018 -218 -1012
rect 76 -977 83 -970
rect 100 -977 107 -970
rect 133 -974 141 -965
rect 187 -974 195 -965
rect -200 -1018 -193 -1012
rect -152 -1018 -144 -1012
rect -134 -1018 -125 -1012
rect 243 -980 250 -973
rect 264 -980 271 -973
rect 375 -977 382 -970
rect 396 -977 403 -970
rect 432 -974 440 -965
rect 486 -974 494 -965
rect 52 -1049 60 -1040
rect 106 -1049 114 -1040
rect -249 -1090 -241 -1081
rect -195 -1090 -187 -1081
rect -166 -1090 -158 -1081
rect -137 -1090 -130 -1081
rect 157 -1062 164 -1055
rect 542 -980 549 -973
rect 563 -980 570 -973
rect 690 -977 697 -970
rect 711 -977 718 -970
rect 747 -974 755 -965
rect 801 -974 809 -965
rect 219 -1052 227 -1043
rect 273 -1052 281 -1043
rect 351 -1049 359 -1040
rect 405 -1049 413 -1040
rect 181 -1062 188 -1055
rect -225 -1121 -218 -1115
rect -202 -1121 -195 -1115
rect -152 -1121 -144 -1115
rect -134 -1121 -125 -1115
rect 80 -1168 87 -1162
rect 101 -1168 108 -1162
rect 456 -1062 463 -1055
rect 857 -980 864 -973
rect 878 -980 885 -973
rect 1019 -971 1026 -964
rect 1040 -971 1047 -964
rect 1076 -968 1084 -959
rect 1130 -968 1138 -959
rect 518 -1052 526 -1043
rect 572 -1052 580 -1043
rect 666 -1049 674 -1040
rect 720 -1049 728 -1040
rect 480 -1062 487 -1055
rect 133 -1134 141 -1125
rect 187 -1134 195 -1125
rect 153 -1168 161 -1162
rect 171 -1168 180 -1162
rect 379 -1168 386 -1162
rect 400 -1168 407 -1162
rect 771 -1062 778 -1055
rect 1186 -974 1193 -967
rect 1207 -974 1214 -967
rect 1334 -971 1341 -964
rect 1355 -971 1362 -964
rect 1391 -968 1399 -959
rect 1445 -968 1453 -959
rect 995 -1043 1003 -1034
rect 1049 -1043 1057 -1034
rect 833 -1052 841 -1043
rect 887 -1052 895 -1043
rect 795 -1062 802 -1055
rect 432 -1134 440 -1125
rect 486 -1134 494 -1125
rect 452 -1168 460 -1162
rect 470 -1168 479 -1162
rect 694 -1168 701 -1162
rect 715 -1168 722 -1162
rect 1100 -1056 1107 -1049
rect 1501 -974 1508 -967
rect 1522 -974 1529 -967
rect 1162 -1046 1170 -1037
rect 1216 -1046 1224 -1037
rect 1310 -1043 1318 -1034
rect 1364 -1043 1372 -1034
rect 1124 -1056 1131 -1049
rect 747 -1134 755 -1125
rect 801 -1134 809 -1125
rect 1023 -1162 1030 -1156
rect 1044 -1162 1051 -1156
rect 767 -1168 775 -1162
rect 785 -1168 794 -1162
rect 1415 -1056 1422 -1049
rect 1477 -1046 1485 -1037
rect 1531 -1046 1539 -1037
rect 1439 -1056 1446 -1049
rect 1076 -1128 1084 -1119
rect 1130 -1128 1138 -1119
rect 1096 -1162 1104 -1156
rect 1114 -1162 1123 -1156
rect 1338 -1162 1345 -1156
rect 1359 -1162 1366 -1156
rect 1391 -1128 1399 -1119
rect 1445 -1128 1453 -1119
rect 1411 -1162 1419 -1156
rect 1429 -1162 1438 -1156
rect -249 -1193 -241 -1184
rect -195 -1193 -187 -1184
rect -166 -1193 -158 -1184
rect -137 -1193 -130 -1184
rect -225 -1221 -218 -1215
rect -200 -1221 -193 -1215
rect -152 -1221 -144 -1215
rect -134 -1221 -125 -1215
rect 831 -1193 837 -1187
rect 857 -1193 863 -1187
rect 884 -1193 890 -1187
rect 903 -1193 909 -1187
rect 56 -1240 64 -1231
rect 110 -1240 118 -1231
rect 139 -1240 147 -1231
rect 168 -1240 175 -1231
rect 355 -1240 363 -1231
rect 409 -1240 417 -1231
rect 438 -1240 446 -1231
rect 467 -1240 474 -1231
rect 670 -1240 678 -1231
rect 724 -1240 732 -1231
rect 753 -1240 761 -1231
rect 782 -1240 789 -1231
rect 157 -1276 164 -1269
rect 178 -1276 185 -1269
rect 1475 -1187 1481 -1181
rect 1501 -1187 1507 -1181
rect 1528 -1187 1534 -1181
rect 1547 -1187 1553 -1181
rect 999 -1234 1007 -1225
rect 1053 -1234 1061 -1225
rect 1082 -1234 1090 -1225
rect 1111 -1234 1118 -1225
rect 1314 -1234 1322 -1225
rect 1368 -1234 1376 -1225
rect 1397 -1234 1405 -1225
rect 1426 -1234 1433 -1225
rect 821 -1259 826 -1254
rect 841 -1259 847 -1254
rect 867 -1259 872 -1254
rect 890 -1259 896 -1254
rect 916 -1259 921 -1254
rect 1465 -1253 1470 -1248
rect 1485 -1253 1491 -1248
rect 1511 -1253 1516 -1248
rect 1534 -1253 1540 -1248
rect 1560 -1253 1565 -1248
rect -249 -1293 -241 -1284
rect -195 -1293 -187 -1284
rect -166 -1293 -158 -1284
rect -137 -1293 -130 -1284
rect -225 -1328 -218 -1322
rect -200 -1328 -193 -1322
rect -152 -1328 -144 -1322
rect -134 -1328 -125 -1322
rect 76 -1351 83 -1344
rect 488 -1309 495 -1302
rect 509 -1309 516 -1302
rect 803 -1309 810 -1302
rect 824 -1309 831 -1302
rect 101 -1351 108 -1344
rect 133 -1348 141 -1339
rect 187 -1348 195 -1339
rect -249 -1400 -241 -1391
rect -195 -1400 -187 -1391
rect -166 -1400 -158 -1391
rect -137 -1400 -130 -1391
rect -225 -1428 -218 -1422
rect 243 -1354 250 -1347
rect 264 -1354 271 -1347
rect -201 -1428 -195 -1422
rect -152 -1428 -144 -1422
rect -134 -1428 -125 -1422
rect 52 -1423 60 -1414
rect 106 -1423 114 -1414
rect 157 -1436 164 -1429
rect 407 -1384 414 -1377
rect 428 -1384 435 -1377
rect 464 -1381 472 -1372
rect 518 -1381 526 -1372
rect 219 -1426 227 -1417
rect 273 -1426 281 -1417
rect 181 -1436 188 -1429
rect -249 -1500 -241 -1491
rect -195 -1500 -187 -1491
rect -166 -1500 -158 -1491
rect -137 -1500 -130 -1491
rect 80 -1542 87 -1536
rect 101 -1542 108 -1536
rect 574 -1387 581 -1380
rect 595 -1387 602 -1380
rect 722 -1384 729 -1377
rect 743 -1384 750 -1377
rect 779 -1381 787 -1372
rect 833 -1381 841 -1372
rect 383 -1456 391 -1447
rect 437 -1456 445 -1447
rect 133 -1508 141 -1499
rect 187 -1508 195 -1499
rect 488 -1469 495 -1462
rect 889 -1387 896 -1380
rect 910 -1387 917 -1380
rect 550 -1459 558 -1450
rect 604 -1459 612 -1450
rect 698 -1456 706 -1447
rect 752 -1456 760 -1447
rect 512 -1469 519 -1462
rect 153 -1542 161 -1536
rect 171 -1542 180 -1536
rect 411 -1575 418 -1569
rect 432 -1575 439 -1569
rect 803 -1469 810 -1462
rect 865 -1459 873 -1450
rect 919 -1459 927 -1450
rect 827 -1469 834 -1462
rect 464 -1541 472 -1532
rect 518 -1541 526 -1532
rect 484 -1575 492 -1569
rect 502 -1575 511 -1569
rect 726 -1575 733 -1569
rect 747 -1575 754 -1569
rect 779 -1541 787 -1532
rect 833 -1541 841 -1532
rect 799 -1575 807 -1569
rect 817 -1575 826 -1569
rect 56 -1614 64 -1605
rect 110 -1614 118 -1605
rect 139 -1614 147 -1605
rect 168 -1614 175 -1605
rect 863 -1600 869 -1594
rect 889 -1600 895 -1594
rect 916 -1600 922 -1594
rect 935 -1600 941 -1594
rect 157 -1652 164 -1645
rect 178 -1652 185 -1645
rect 387 -1647 395 -1638
rect 441 -1647 449 -1638
rect 470 -1647 478 -1638
rect 499 -1647 506 -1638
rect 702 -1647 710 -1638
rect 756 -1647 764 -1638
rect 785 -1647 793 -1638
rect 814 -1647 821 -1638
rect 76 -1727 83 -1720
rect 853 -1666 858 -1661
rect 873 -1666 879 -1661
rect 899 -1666 904 -1661
rect 922 -1666 928 -1661
rect 948 -1666 953 -1661
rect 101 -1727 108 -1720
rect 133 -1724 141 -1715
rect 187 -1724 195 -1715
rect 243 -1730 250 -1723
rect 264 -1730 271 -1723
rect 52 -1799 60 -1790
rect 106 -1799 114 -1790
rect 157 -1812 164 -1805
rect 219 -1802 227 -1793
rect 273 -1802 281 -1793
rect 181 -1812 188 -1805
rect 80 -1918 87 -1912
rect 101 -1918 108 -1912
rect 133 -1884 141 -1875
rect 187 -1884 195 -1875
rect 153 -1918 161 -1912
rect 171 -1918 180 -1912
rect 56 -1990 64 -1981
rect 110 -1990 118 -1981
rect 139 -1990 147 -1981
rect 168 -1990 175 -1981
<< pdcontact >>
rect 138 352 145 360
rect 160 352 167 360
rect 187 352 194 360
rect 425 352 432 360
rect 447 352 454 360
rect 474 352 481 360
rect 57 277 64 285
rect 79 277 86 285
rect 106 277 113 285
rect 224 274 231 282
rect 246 274 253 282
rect 273 274 280 282
rect 344 277 351 285
rect 366 277 373 285
rect 393 277 400 285
rect 511 274 518 282
rect 533 274 540 282
rect 560 274 567 282
rect 138 192 145 200
rect 160 192 167 200
rect 187 192 194 200
rect 425 192 432 200
rect 447 192 454 200
rect 474 192 481 200
rect -243 98 -236 106
rect -221 98 -214 106
rect -194 98 -187 106
rect -158 98 -151 106
rect -136 98 -129 106
rect 61 86 68 94
rect 83 86 90 94
rect 110 86 117 94
rect 146 86 153 94
rect 168 86 175 94
rect 348 86 355 94
rect 370 86 377 94
rect 397 86 404 94
rect 433 86 440 94
rect 455 86 462 94
rect 495 80 500 89
rect 541 80 546 89
rect 568 80 573 89
rect 589 80 594 89
rect 500 20 506 26
rect 531 20 537 26
rect 553 20 559 26
rect 572 20 578 26
rect -243 -2 -236 6
rect -221 -2 -214 6
rect -194 -2 -187 6
rect -158 -2 -151 6
rect -136 -2 -129 6
rect 138 -51 145 -43
rect 160 -51 167 -43
rect 187 -51 194 -43
rect 425 -51 432 -43
rect 447 -51 454 -43
rect 474 -51 481 -43
rect 770 -50 777 -42
rect 792 -50 799 -42
rect 819 -50 826 -42
rect 1085 -50 1092 -42
rect 1107 -50 1114 -42
rect 1134 -50 1141 -42
rect -243 -109 -236 -101
rect -221 -109 -214 -101
rect -194 -109 -187 -101
rect -158 -109 -151 -101
rect -136 -109 -129 -101
rect 57 -126 64 -118
rect 79 -126 86 -118
rect 106 -126 113 -118
rect 224 -129 231 -121
rect 246 -129 253 -121
rect 273 -129 280 -121
rect 344 -126 351 -118
rect 366 -126 373 -118
rect 393 -126 400 -118
rect -243 -209 -236 -201
rect -221 -209 -214 -201
rect -194 -209 -187 -201
rect -158 -209 -151 -201
rect -136 -209 -129 -201
rect 511 -129 518 -121
rect 533 -129 540 -121
rect 560 -129 567 -121
rect 689 -125 696 -117
rect 711 -125 718 -117
rect 738 -125 745 -117
rect 138 -211 145 -203
rect 160 -211 167 -203
rect 187 -211 194 -203
rect 856 -128 863 -120
rect 878 -128 885 -120
rect 905 -128 912 -120
rect 1004 -125 1011 -117
rect 1026 -125 1033 -117
rect 1053 -125 1060 -117
rect 425 -211 432 -203
rect 447 -211 454 -203
rect 474 -211 481 -203
rect 1171 -128 1178 -120
rect 1193 -128 1200 -120
rect 1220 -128 1227 -120
rect 770 -210 777 -202
rect 792 -210 799 -202
rect 819 -210 826 -202
rect -243 -312 -236 -304
rect -221 -312 -214 -304
rect -194 -312 -187 -304
rect -158 -312 -151 -304
rect -136 -312 -129 -304
rect 61 -317 68 -309
rect 83 -317 90 -309
rect 110 -317 117 -309
rect 146 -317 153 -309
rect 168 -317 175 -309
rect 348 -317 355 -309
rect 370 -317 377 -309
rect 397 -317 404 -309
rect 433 -317 440 -309
rect 455 -317 462 -309
rect 1085 -210 1092 -202
rect 1107 -210 1114 -202
rect 1134 -210 1141 -202
rect 495 -323 500 -314
rect 541 -323 546 -314
rect 568 -323 573 -314
rect 589 -323 594 -314
rect 693 -316 700 -308
rect 715 -316 722 -308
rect 742 -316 749 -308
rect 778 -316 785 -308
rect 800 -316 807 -308
rect 1008 -316 1015 -308
rect 1030 -316 1037 -308
rect 1057 -316 1064 -308
rect 1093 -316 1100 -308
rect 1115 -316 1122 -308
rect 1155 -322 1160 -313
rect 1201 -322 1206 -313
rect 1228 -322 1233 -313
rect 1249 -322 1254 -313
rect 500 -383 506 -377
rect 531 -383 537 -377
rect 553 -383 559 -377
rect 572 -383 578 -377
rect 1160 -382 1166 -376
rect 1191 -382 1197 -376
rect 1213 -382 1219 -376
rect 1232 -382 1238 -376
rect -243 -412 -236 -404
rect -221 -412 -214 -404
rect -194 -412 -187 -404
rect -158 -412 -151 -404
rect -136 -412 -129 -404
rect 138 -467 145 -459
rect 160 -467 167 -459
rect 187 -467 194 -459
rect 425 -467 432 -459
rect 447 -467 454 -459
rect 474 -467 481 -459
rect 771 -467 778 -459
rect 793 -467 800 -459
rect 820 -467 827 -459
rect 1053 -467 1060 -459
rect 1075 -467 1082 -459
rect 1102 -467 1109 -459
rect 1380 -462 1387 -454
rect 1402 -462 1409 -454
rect 1429 -462 1436 -454
rect -243 -519 -236 -511
rect -221 -519 -214 -511
rect -194 -519 -187 -511
rect -158 -519 -151 -511
rect -136 -519 -129 -511
rect 57 -542 64 -534
rect 79 -542 86 -534
rect 106 -542 113 -534
rect 224 -545 231 -537
rect 246 -545 253 -537
rect 273 -545 280 -537
rect 344 -542 351 -534
rect 366 -542 373 -534
rect 393 -542 400 -534
rect -243 -619 -236 -611
rect -221 -619 -214 -611
rect -194 -619 -187 -611
rect -158 -619 -151 -611
rect -136 -619 -129 -611
rect 511 -545 518 -537
rect 533 -545 540 -537
rect 560 -545 567 -537
rect 690 -542 697 -534
rect 712 -542 719 -534
rect 739 -542 746 -534
rect 138 -627 145 -619
rect 160 -627 167 -619
rect 187 -627 194 -619
rect 857 -545 864 -537
rect 879 -545 886 -537
rect 906 -545 913 -537
rect 972 -542 979 -534
rect 994 -542 1001 -534
rect 1021 -542 1028 -534
rect 425 -627 432 -619
rect 447 -627 454 -619
rect 474 -627 481 -619
rect 1299 -537 1306 -529
rect 1321 -537 1328 -529
rect 1348 -537 1355 -529
rect 1139 -545 1146 -537
rect 1161 -545 1168 -537
rect 1188 -545 1195 -537
rect 771 -627 778 -619
rect 793 -627 800 -619
rect 820 -627 827 -619
rect -244 -734 -237 -726
rect -222 -734 -215 -726
rect -195 -734 -188 -726
rect -159 -734 -152 -726
rect -137 -734 -130 -726
rect 61 -733 68 -725
rect 83 -733 90 -725
rect 110 -733 117 -725
rect 146 -733 153 -725
rect 168 -733 175 -725
rect 348 -733 355 -725
rect 370 -733 377 -725
rect 397 -733 404 -725
rect 433 -733 440 -725
rect 455 -733 462 -725
rect 1466 -540 1473 -532
rect 1488 -540 1495 -532
rect 1515 -540 1522 -532
rect 1053 -627 1060 -619
rect 1075 -627 1082 -619
rect 1102 -627 1109 -619
rect 1380 -622 1387 -614
rect 1402 -622 1409 -614
rect 1429 -622 1436 -614
rect 495 -739 500 -730
rect 541 -739 546 -730
rect 568 -739 573 -730
rect 589 -739 594 -730
rect 694 -733 701 -725
rect 716 -733 723 -725
rect 743 -733 750 -725
rect 779 -733 786 -725
rect 801 -733 808 -725
rect 976 -733 983 -725
rect 998 -733 1005 -725
rect 1025 -733 1032 -725
rect 1061 -733 1068 -725
rect 1083 -733 1090 -725
rect 1303 -728 1310 -720
rect 1325 -728 1332 -720
rect 1352 -728 1359 -720
rect 1388 -728 1395 -720
rect 1410 -728 1417 -720
rect 1123 -739 1128 -730
rect 1169 -739 1174 -730
rect 1196 -739 1201 -730
rect 1217 -739 1222 -730
rect 500 -799 506 -793
rect 531 -799 537 -793
rect 553 -799 559 -793
rect 572 -799 578 -793
rect 1128 -799 1134 -793
rect 1159 -799 1165 -793
rect 1181 -799 1187 -793
rect 1200 -799 1206 -793
rect -244 -834 -237 -826
rect -222 -834 -215 -826
rect -195 -834 -188 -826
rect -159 -834 -152 -826
rect -137 -834 -130 -826
rect 138 -925 145 -917
rect 160 -925 167 -917
rect 187 -925 194 -917
rect 437 -925 444 -917
rect 459 -925 466 -917
rect 486 -925 493 -917
rect 752 -925 759 -917
rect 774 -925 781 -917
rect 801 -925 808 -917
rect 1081 -919 1088 -911
rect 1103 -919 1110 -911
rect 1130 -919 1137 -911
rect 1396 -919 1403 -911
rect 1418 -919 1425 -911
rect 1445 -919 1452 -911
rect -244 -941 -237 -933
rect -222 -941 -215 -933
rect -195 -941 -188 -933
rect -159 -941 -152 -933
rect -137 -941 -130 -933
rect 57 -1000 64 -992
rect 79 -1000 86 -992
rect 106 -1000 113 -992
rect -244 -1041 -237 -1033
rect -222 -1041 -215 -1033
rect -195 -1041 -188 -1033
rect -159 -1041 -152 -1033
rect -137 -1041 -130 -1033
rect 224 -1003 231 -995
rect 246 -1003 253 -995
rect 273 -1003 280 -995
rect 356 -1000 363 -992
rect 378 -1000 385 -992
rect 405 -1000 412 -992
rect 523 -1003 530 -995
rect 545 -1003 552 -995
rect 572 -1003 579 -995
rect 671 -1000 678 -992
rect 693 -1000 700 -992
rect 720 -1000 727 -992
rect 138 -1085 145 -1077
rect 160 -1085 167 -1077
rect 187 -1085 194 -1077
rect -244 -1144 -237 -1136
rect -222 -1144 -215 -1136
rect -195 -1144 -188 -1136
rect -159 -1144 -152 -1136
rect -137 -1144 -130 -1136
rect 1000 -994 1007 -986
rect 1022 -994 1029 -986
rect 1049 -994 1056 -986
rect 838 -1003 845 -995
rect 860 -1003 867 -995
rect 887 -1003 894 -995
rect 437 -1085 444 -1077
rect 459 -1085 466 -1077
rect 486 -1085 493 -1077
rect 1167 -997 1174 -989
rect 1189 -997 1196 -989
rect 1216 -997 1223 -989
rect 1315 -994 1322 -986
rect 1337 -994 1344 -986
rect 1364 -994 1371 -986
rect 752 -1085 759 -1077
rect 774 -1085 781 -1077
rect 801 -1085 808 -1077
rect 1482 -997 1489 -989
rect 1504 -997 1511 -989
rect 1531 -997 1538 -989
rect 1081 -1079 1088 -1071
rect 1103 -1079 1110 -1071
rect 1130 -1079 1137 -1071
rect 1396 -1079 1403 -1071
rect 1418 -1079 1425 -1071
rect 1445 -1079 1452 -1071
rect 61 -1191 68 -1183
rect 83 -1191 90 -1183
rect 110 -1191 117 -1183
rect 146 -1191 153 -1183
rect 168 -1191 175 -1183
rect 360 -1191 367 -1183
rect 382 -1191 389 -1183
rect 409 -1191 416 -1183
rect 445 -1191 452 -1183
rect 467 -1191 474 -1183
rect 675 -1191 682 -1183
rect 697 -1191 704 -1183
rect 724 -1191 731 -1183
rect 760 -1191 767 -1183
rect 782 -1191 789 -1183
rect 1004 -1185 1011 -1177
rect 1026 -1185 1033 -1177
rect 1053 -1185 1060 -1177
rect 1089 -1185 1096 -1177
rect 1111 -1185 1118 -1177
rect 1319 -1185 1326 -1177
rect 1341 -1185 1348 -1177
rect 1368 -1185 1375 -1177
rect 1404 -1185 1411 -1177
rect 1426 -1185 1433 -1177
rect 822 -1217 827 -1208
rect 868 -1217 873 -1208
rect 895 -1217 900 -1208
rect 916 -1217 921 -1208
rect -244 -1244 -237 -1236
rect -222 -1244 -215 -1236
rect -195 -1244 -188 -1236
rect -159 -1244 -152 -1236
rect -137 -1244 -130 -1236
rect 1466 -1211 1471 -1202
rect 1512 -1211 1517 -1202
rect 1539 -1211 1544 -1202
rect 1560 -1211 1565 -1202
rect 827 -1277 833 -1271
rect 858 -1277 864 -1271
rect 880 -1277 886 -1271
rect 899 -1277 905 -1271
rect 1471 -1271 1477 -1265
rect 1502 -1271 1508 -1265
rect 1524 -1271 1530 -1265
rect 1543 -1271 1549 -1265
rect 138 -1299 145 -1291
rect 160 -1299 167 -1291
rect 187 -1299 194 -1291
rect -244 -1351 -237 -1343
rect -222 -1351 -215 -1343
rect -195 -1351 -188 -1343
rect -159 -1351 -152 -1343
rect -137 -1351 -130 -1343
rect 57 -1374 64 -1366
rect 79 -1374 86 -1366
rect 106 -1374 113 -1366
rect 469 -1332 476 -1324
rect 491 -1332 498 -1324
rect 518 -1332 525 -1324
rect 784 -1332 791 -1324
rect 806 -1332 813 -1324
rect 833 -1332 840 -1324
rect 224 -1377 231 -1369
rect 246 -1377 253 -1369
rect 273 -1377 280 -1369
rect -244 -1451 -237 -1443
rect -222 -1451 -215 -1443
rect -195 -1451 -188 -1443
rect -159 -1451 -152 -1443
rect -137 -1451 -130 -1443
rect 388 -1407 395 -1399
rect 410 -1407 417 -1399
rect 437 -1407 444 -1399
rect 138 -1459 145 -1451
rect 160 -1459 167 -1451
rect 187 -1459 194 -1451
rect 555 -1410 562 -1402
rect 577 -1410 584 -1402
rect 604 -1410 611 -1402
rect 703 -1407 710 -1399
rect 725 -1407 732 -1399
rect 752 -1407 759 -1399
rect 870 -1410 877 -1402
rect 892 -1410 899 -1402
rect 919 -1410 926 -1402
rect 469 -1492 476 -1484
rect 491 -1492 498 -1484
rect 518 -1492 525 -1484
rect 61 -1565 68 -1557
rect 83 -1565 90 -1557
rect 110 -1565 117 -1557
rect 146 -1565 153 -1557
rect 168 -1565 175 -1557
rect 784 -1492 791 -1484
rect 806 -1492 813 -1484
rect 833 -1492 840 -1484
rect 392 -1598 399 -1590
rect 414 -1598 421 -1590
rect 441 -1598 448 -1590
rect 477 -1598 484 -1590
rect 499 -1598 506 -1590
rect 707 -1598 714 -1590
rect 729 -1598 736 -1590
rect 756 -1598 763 -1590
rect 792 -1598 799 -1590
rect 814 -1598 821 -1590
rect 854 -1624 859 -1615
rect 900 -1624 905 -1615
rect 927 -1624 932 -1615
rect 948 -1624 953 -1615
rect 138 -1675 145 -1667
rect 160 -1675 167 -1667
rect 187 -1675 194 -1667
rect 859 -1684 865 -1678
rect 890 -1684 896 -1678
rect 912 -1684 918 -1678
rect 931 -1684 937 -1678
rect 57 -1750 64 -1742
rect 79 -1750 86 -1742
rect 106 -1750 113 -1742
rect 224 -1753 231 -1745
rect 246 -1753 253 -1745
rect 273 -1753 280 -1745
rect 138 -1835 145 -1827
rect 160 -1835 167 -1827
rect 187 -1835 194 -1827
rect 61 -1941 68 -1933
rect 83 -1941 90 -1933
rect 110 -1941 117 -1933
rect 146 -1941 153 -1933
rect 168 -1941 175 -1933
<< psubstratepcontact >>
rect 145 286 153 294
rect 432 286 440 294
rect 64 211 72 219
rect 231 208 239 216
rect 351 211 359 219
rect 518 208 526 216
rect 145 126 153 134
rect 173 126 181 134
rect 432 126 440 134
rect 460 126 468 134
rect -236 32 -228 40
rect -200 32 -192 40
rect -157 32 -148 40
rect -138 32 -129 40
rect 68 20 76 28
rect 105 20 113 28
rect 147 20 156 28
rect 166 20 175 28
rect 355 20 363 28
rect 383 20 391 28
rect 434 20 443 28
rect 453 20 462 28
rect -236 -68 -228 -60
rect -200 -68 -192 -60
rect -157 -68 -148 -60
rect -138 -68 -129 -60
rect 145 -117 153 -109
rect -236 -175 -228 -167
rect 432 -117 440 -109
rect -200 -175 -192 -167
rect -157 -175 -148 -167
rect -138 -175 -129 -167
rect 64 -192 72 -184
rect 777 -116 785 -108
rect 231 -195 239 -187
rect -236 -275 -228 -267
rect -200 -275 -192 -267
rect -157 -275 -148 -267
rect -138 -275 -129 -267
rect 351 -192 359 -184
rect 1092 -116 1100 -108
rect 518 -195 526 -187
rect 145 -277 153 -269
rect 173 -277 181 -269
rect 696 -191 704 -183
rect 863 -194 871 -186
rect 432 -277 440 -269
rect 460 -277 468 -269
rect 1011 -191 1019 -183
rect 1178 -194 1186 -186
rect 777 -276 785 -268
rect 805 -276 813 -268
rect 1092 -276 1100 -268
rect 1120 -276 1128 -268
rect -236 -378 -228 -370
rect -200 -378 -192 -370
rect -157 -378 -148 -370
rect -138 -378 -129 -370
rect 68 -383 76 -375
rect 105 -383 113 -375
rect 147 -383 156 -375
rect 166 -383 175 -375
rect 355 -383 363 -375
rect 391 -383 399 -375
rect 434 -383 443 -375
rect 453 -383 462 -375
rect 700 -382 708 -374
rect 737 -382 745 -374
rect 779 -382 788 -374
rect 798 -382 807 -374
rect 1015 -382 1023 -374
rect 1051 -382 1059 -374
rect 1094 -382 1103 -374
rect 1113 -382 1122 -374
rect -236 -478 -228 -470
rect -200 -478 -192 -470
rect -157 -478 -148 -470
rect -138 -478 -129 -470
rect 145 -533 153 -525
rect -236 -585 -228 -577
rect -200 -585 -192 -577
rect -157 -585 -148 -577
rect -138 -585 -129 -577
rect 432 -533 440 -525
rect 64 -608 72 -600
rect 778 -533 786 -525
rect 231 -611 239 -603
rect -236 -685 -228 -677
rect -200 -685 -192 -677
rect -157 -685 -148 -677
rect -138 -685 -129 -677
rect 351 -608 359 -600
rect 1060 -533 1068 -525
rect 518 -611 526 -603
rect 145 -693 153 -685
rect 173 -693 181 -685
rect 697 -608 705 -600
rect 1387 -528 1395 -520
rect 864 -611 872 -603
rect 432 -693 440 -685
rect 460 -693 468 -685
rect 979 -608 987 -600
rect 1146 -611 1154 -603
rect 778 -693 786 -685
rect 806 -693 814 -685
rect 1306 -603 1314 -595
rect 1473 -606 1481 -598
rect 1060 -693 1068 -685
rect 1088 -693 1096 -685
rect 1387 -688 1395 -680
rect 1415 -688 1423 -680
rect -237 -800 -229 -792
rect -201 -800 -193 -792
rect -158 -800 -149 -792
rect -139 -800 -130 -792
rect 68 -799 76 -791
rect 105 -799 113 -791
rect 147 -799 156 -791
rect 166 -799 175 -791
rect 355 -799 363 -791
rect 391 -799 399 -791
rect 434 -799 443 -791
rect 453 -799 462 -791
rect 701 -799 709 -791
rect 738 -799 746 -791
rect 780 -799 789 -791
rect 799 -799 808 -791
rect 983 -799 991 -791
rect 1019 -799 1027 -791
rect 1062 -799 1071 -791
rect 1081 -799 1090 -791
rect 1310 -794 1318 -786
rect 1348 -794 1356 -786
rect 1389 -794 1398 -786
rect 1408 -794 1417 -786
rect -237 -900 -229 -892
rect -201 -900 -193 -892
rect -158 -900 -149 -892
rect -139 -900 -130 -892
rect -237 -1007 -229 -999
rect 145 -991 153 -983
rect -201 -1007 -193 -999
rect -158 -1007 -149 -999
rect -139 -1007 -130 -999
rect 444 -991 452 -983
rect 64 -1066 72 -1058
rect 759 -991 767 -983
rect 231 -1069 239 -1061
rect -237 -1107 -229 -1099
rect -201 -1107 -193 -1099
rect -158 -1107 -149 -1099
rect -139 -1107 -130 -1099
rect 363 -1066 371 -1058
rect 1088 -985 1096 -977
rect 530 -1069 538 -1061
rect 145 -1151 153 -1143
rect 173 -1151 181 -1143
rect 678 -1066 686 -1058
rect 1403 -985 1411 -977
rect 845 -1069 853 -1061
rect 444 -1151 452 -1143
rect 472 -1151 480 -1143
rect 1007 -1060 1015 -1052
rect 1174 -1063 1182 -1055
rect 759 -1151 767 -1143
rect 787 -1151 795 -1143
rect 1322 -1060 1330 -1052
rect 1489 -1063 1497 -1055
rect 1088 -1145 1096 -1137
rect 1116 -1145 1124 -1137
rect 1403 -1145 1411 -1137
rect 1431 -1145 1439 -1137
rect -237 -1210 -229 -1202
rect -201 -1210 -193 -1202
rect -158 -1210 -149 -1202
rect -139 -1210 -130 -1202
rect 68 -1257 76 -1249
rect 96 -1257 104 -1249
rect 147 -1257 156 -1249
rect 166 -1257 175 -1249
rect 367 -1257 375 -1249
rect 404 -1257 412 -1249
rect 446 -1257 455 -1249
rect 465 -1257 474 -1249
rect 682 -1257 690 -1249
rect 719 -1257 727 -1249
rect 761 -1257 770 -1249
rect 780 -1257 789 -1249
rect 1011 -1251 1019 -1243
rect 1048 -1251 1056 -1243
rect 1090 -1251 1099 -1243
rect 1109 -1251 1118 -1243
rect 1326 -1251 1334 -1243
rect 1362 -1251 1370 -1243
rect 1405 -1251 1414 -1243
rect 1424 -1251 1433 -1243
rect -237 -1310 -229 -1302
rect -201 -1310 -193 -1302
rect -158 -1310 -149 -1302
rect -139 -1310 -130 -1302
rect 145 -1365 153 -1357
rect -237 -1417 -229 -1409
rect -201 -1417 -193 -1409
rect -158 -1417 -149 -1409
rect -139 -1417 -130 -1409
rect 64 -1440 72 -1432
rect 476 -1398 484 -1390
rect 231 -1443 239 -1435
rect -237 -1517 -229 -1509
rect -201 -1517 -193 -1509
rect -158 -1517 -149 -1509
rect -139 -1517 -130 -1509
rect 791 -1398 799 -1390
rect 395 -1473 403 -1465
rect 562 -1476 570 -1468
rect 145 -1525 153 -1517
rect 173 -1525 181 -1517
rect 710 -1473 718 -1465
rect 877 -1476 885 -1468
rect 476 -1558 484 -1550
rect 504 -1558 512 -1550
rect 791 -1558 799 -1550
rect 819 -1558 827 -1550
rect 68 -1631 76 -1623
rect 96 -1631 104 -1623
rect 147 -1631 156 -1623
rect 166 -1631 175 -1623
rect 399 -1664 407 -1656
rect 436 -1664 444 -1656
rect 478 -1664 487 -1656
rect 497 -1664 506 -1656
rect 714 -1664 722 -1656
rect 750 -1664 758 -1656
rect 793 -1664 802 -1656
rect 812 -1664 821 -1656
rect 145 -1741 153 -1733
rect 64 -1816 72 -1808
rect 231 -1819 239 -1811
rect 145 -1901 153 -1893
rect 173 -1901 181 -1893
rect 68 -2007 76 -1999
rect 96 -2007 104 -1999
rect 147 -2007 156 -1999
rect 166 -2007 175 -1999
<< polysilicon >>
rect 147 360 152 368
rect 175 360 180 368
rect 434 360 439 368
rect 462 360 467 368
rect 147 335 152 352
rect 66 330 70 335
rect 141 330 152 335
rect 66 285 71 330
rect 147 312 152 330
rect 175 312 180 352
rect 195 328 200 336
rect 147 300 152 303
rect 94 285 99 293
rect 66 252 71 277
rect 47 245 71 252
rect 66 237 71 245
rect 94 237 99 277
rect 175 261 180 303
rect 233 282 238 328
rect 353 330 357 335
rect 261 282 266 290
rect 353 285 358 330
rect 381 285 386 343
rect 434 335 439 352
rect 428 330 439 335
rect 434 312 439 330
rect 462 312 467 352
rect 482 328 487 336
rect 434 300 439 303
rect 114 253 180 261
rect 66 225 71 228
rect 94 180 99 228
rect 147 200 152 208
rect 175 200 180 253
rect 233 234 238 274
rect 261 234 266 274
rect 281 252 334 258
rect 353 252 358 277
rect 281 250 326 252
rect 334 245 358 252
rect 353 237 358 245
rect 381 237 386 277
rect 462 261 467 303
rect 520 282 525 328
rect 548 282 553 290
rect 401 253 467 261
rect 353 225 358 228
rect 233 222 238 225
rect 94 163 98 180
rect 94 159 115 163
rect -234 106 -229 114
rect -206 106 -201 114
rect -149 106 -144 114
rect 111 107 115 159
rect 147 152 152 192
rect 175 152 180 192
rect 261 176 266 225
rect 195 168 266 176
rect 381 180 386 228
rect 434 200 439 208
rect 462 200 467 253
rect 520 234 525 274
rect 548 234 553 274
rect 568 250 576 258
rect 520 222 525 225
rect 381 163 385 180
rect 381 159 402 163
rect 147 140 152 143
rect 175 140 180 143
rect 398 107 402 159
rect 434 152 439 192
rect 462 152 467 192
rect 548 176 553 225
rect 482 168 553 176
rect 434 140 439 143
rect 462 140 467 143
rect 478 113 527 118
rect 98 102 115 107
rect 385 102 402 107
rect -234 74 -229 98
rect -280 68 -229 74
rect -234 58 -229 68
rect -206 58 -201 98
rect -149 82 -144 98
rect 70 94 75 102
rect 98 94 103 102
rect 155 94 160 102
rect 357 94 362 102
rect 385 94 390 102
rect 442 94 447 102
rect -186 74 -144 82
rect -149 58 -144 74
rect 70 63 75 86
rect 47 56 75 63
rect -234 46 -229 49
rect -234 6 -229 14
rect -206 6 -201 49
rect -149 45 -144 49
rect 70 46 75 56
rect 98 46 103 86
rect 155 70 160 86
rect 118 62 160 70
rect 357 63 362 86
rect 155 46 160 62
rect 334 56 362 63
rect 357 46 362 56
rect 385 46 390 86
rect 442 70 447 86
rect 478 71 482 113
rect 521 101 527 113
rect 521 96 534 101
rect 503 89 507 92
rect 530 89 534 96
rect 578 89 583 92
rect 405 62 447 70
rect 467 64 482 71
rect 503 62 507 80
rect 442 46 447 62
rect 504 55 507 62
rect 503 43 507 55
rect 530 43 534 80
rect 578 60 583 80
rect 551 55 583 60
rect 578 43 583 55
rect 70 34 75 37
rect -149 6 -144 14
rect 98 7 103 37
rect 155 33 160 37
rect 357 34 362 37
rect 385 34 390 37
rect 442 33 447 37
rect 503 35 507 38
rect 530 34 534 38
rect 578 34 583 38
rect -234 -29 -229 -2
rect -271 -35 -229 -29
rect -234 -42 -229 -35
rect -206 -42 -201 -2
rect -149 -18 -144 -2
rect -186 -26 -144 -18
rect -149 -42 -144 -26
rect 147 -43 152 -35
rect 175 -43 180 -35
rect 434 -43 439 -35
rect 462 -43 467 -35
rect 779 -42 784 -34
rect 807 -42 812 -34
rect 1094 -42 1099 -34
rect 1122 -42 1127 -34
rect -234 -54 -229 -51
rect -234 -101 -229 -93
rect -206 -101 -201 -51
rect -149 -55 -144 -51
rect 147 -68 152 -51
rect 66 -73 70 -68
rect 141 -73 152 -68
rect -149 -101 -144 -93
rect -234 -131 -229 -109
rect -262 -137 -229 -131
rect -234 -149 -229 -137
rect -206 -149 -201 -109
rect -149 -125 -144 -109
rect 66 -118 71 -73
rect 147 -91 152 -73
rect 175 -91 180 -51
rect 195 -75 200 -67
rect 434 -68 439 -51
rect 147 -103 152 -100
rect 94 -118 99 -110
rect -186 -133 -144 -125
rect -149 -149 -144 -133
rect 66 -151 71 -126
rect 47 -158 71 -151
rect -234 -161 -229 -158
rect -234 -201 -229 -193
rect -206 -201 -201 -158
rect -149 -162 -144 -158
rect 66 -166 71 -158
rect 94 -166 99 -126
rect 175 -142 180 -100
rect 233 -121 238 -75
rect 353 -73 357 -68
rect 428 -73 439 -68
rect 261 -121 266 -113
rect 353 -118 358 -73
rect 434 -91 439 -73
rect 462 -91 467 -51
rect 779 -67 784 -50
rect 482 -75 487 -67
rect 434 -103 439 -100
rect 381 -118 386 -110
rect 114 -150 180 -142
rect 66 -178 71 -175
rect -149 -201 -144 -193
rect -234 -231 -229 -209
rect -253 -237 -229 -231
rect -234 -249 -229 -237
rect -206 -249 -201 -209
rect -149 -225 -144 -209
rect -186 -233 -144 -225
rect -149 -249 -144 -233
rect 94 -223 99 -175
rect 147 -203 152 -195
rect 175 -203 180 -150
rect 233 -169 238 -129
rect 261 -169 266 -129
rect 281 -151 334 -145
rect 353 -151 358 -126
rect 281 -153 326 -151
rect 334 -158 358 -151
rect 353 -166 358 -158
rect 381 -166 386 -126
rect 462 -142 467 -100
rect 520 -121 525 -75
rect 698 -72 702 -67
rect 773 -72 784 -67
rect 548 -121 553 -113
rect 698 -117 703 -72
rect 779 -90 784 -72
rect 807 -90 812 -50
rect 827 -74 832 -66
rect 1094 -67 1099 -50
rect 779 -102 784 -99
rect 726 -117 731 -109
rect 401 -150 467 -142
rect 353 -178 358 -175
rect 233 -181 238 -178
rect 94 -240 98 -223
rect 94 -244 115 -240
rect -234 -261 -229 -258
rect -206 -261 -201 -258
rect -149 -262 -144 -258
rect 111 -296 115 -244
rect 147 -251 152 -211
rect 175 -251 180 -211
rect 261 -227 266 -178
rect 195 -235 266 -227
rect 381 -223 386 -175
rect 434 -203 439 -195
rect 462 -203 467 -150
rect 520 -169 525 -129
rect 548 -169 553 -129
rect 568 -153 619 -145
rect 698 -150 703 -125
rect 679 -157 703 -150
rect 698 -165 703 -157
rect 726 -165 731 -125
rect 807 -141 812 -99
rect 865 -120 870 -74
rect 1013 -72 1017 -67
rect 1088 -72 1099 -67
rect 893 -120 898 -112
rect 1013 -117 1018 -72
rect 1094 -90 1099 -72
rect 1122 -90 1127 -50
rect 1142 -74 1147 -66
rect 1094 -102 1099 -99
rect 1041 -117 1046 -109
rect 746 -149 812 -141
rect 698 -177 703 -174
rect 520 -181 525 -178
rect 381 -240 385 -223
rect 381 -244 402 -240
rect 147 -263 152 -260
rect 175 -263 180 -260
rect 398 -296 402 -244
rect 434 -251 439 -211
rect 462 -251 467 -211
rect 548 -227 553 -178
rect 482 -235 553 -227
rect 726 -222 731 -174
rect 779 -202 784 -194
rect 807 -202 812 -149
rect 865 -168 870 -128
rect 893 -168 898 -128
rect 913 -150 994 -144
rect 1013 -150 1018 -125
rect 913 -152 986 -150
rect 994 -157 1018 -150
rect 1013 -165 1018 -157
rect 1041 -165 1046 -125
rect 1122 -141 1127 -99
rect 1180 -120 1185 -74
rect 1208 -120 1213 -112
rect 1061 -149 1127 -141
rect 1013 -177 1018 -174
rect 865 -180 870 -177
rect 726 -239 730 -222
rect 726 -243 747 -239
rect 434 -263 439 -260
rect 462 -263 467 -260
rect 478 -292 527 -289
rect -234 -304 -229 -296
rect -206 -304 -201 -296
rect -149 -304 -144 -296
rect 98 -301 115 -296
rect 385 -301 402 -296
rect 70 -309 75 -301
rect 98 -309 103 -301
rect 155 -309 160 -301
rect 357 -309 362 -301
rect 385 -309 390 -301
rect 442 -309 447 -301
rect -234 -328 -229 -312
rect -280 -334 -229 -328
rect -234 -352 -229 -334
rect -206 -352 -201 -312
rect -149 -328 -144 -312
rect -186 -336 -144 -328
rect -149 -352 -144 -336
rect 70 -340 75 -317
rect 47 -347 75 -340
rect 70 -357 75 -347
rect 98 -357 103 -317
rect 155 -333 160 -317
rect 118 -341 160 -333
rect 357 -340 362 -317
rect 155 -357 160 -341
rect 334 -347 362 -340
rect 357 -357 362 -347
rect 385 -357 390 -317
rect 442 -333 447 -317
rect 478 -332 482 -292
rect 523 -302 527 -292
rect 743 -295 747 -243
rect 779 -250 784 -210
rect 807 -250 812 -210
rect 893 -226 898 -177
rect 827 -234 898 -226
rect 1041 -222 1046 -174
rect 1094 -202 1099 -194
rect 1122 -202 1127 -149
rect 1180 -168 1185 -128
rect 1208 -168 1213 -128
rect 1228 -152 1236 -144
rect 1180 -180 1185 -177
rect 1041 -239 1045 -222
rect 1041 -243 1062 -239
rect 779 -262 784 -259
rect 807 -262 812 -259
rect 1058 -295 1062 -243
rect 1094 -250 1099 -210
rect 1122 -250 1127 -210
rect 1208 -226 1213 -177
rect 1142 -234 1213 -226
rect 1094 -262 1099 -259
rect 1122 -262 1127 -259
rect 1137 -291 1187 -284
rect 730 -300 747 -295
rect 1045 -300 1062 -295
rect 523 -305 534 -302
rect 503 -314 507 -311
rect 530 -314 534 -305
rect 702 -308 707 -300
rect 730 -308 735 -300
rect 787 -308 792 -300
rect 1017 -308 1022 -300
rect 1045 -308 1050 -300
rect 1102 -308 1107 -300
rect 578 -314 583 -311
rect 405 -341 447 -333
rect 467 -339 482 -332
rect 503 -341 507 -323
rect 442 -357 447 -341
rect 504 -348 507 -341
rect -234 -364 -229 -361
rect -234 -404 -229 -396
rect -206 -404 -201 -361
rect -149 -365 -144 -361
rect 503 -360 507 -348
rect 530 -360 534 -323
rect 578 -343 583 -323
rect 702 -339 707 -316
rect 551 -348 583 -343
rect 679 -346 707 -339
rect 578 -360 583 -348
rect 702 -356 707 -346
rect 730 -356 735 -316
rect 787 -332 792 -316
rect 750 -340 792 -332
rect 1017 -339 1022 -316
rect 787 -356 792 -340
rect 994 -346 1022 -339
rect 1017 -356 1022 -346
rect 1045 -356 1050 -316
rect 1102 -332 1107 -316
rect 1137 -331 1141 -291
rect 1181 -301 1187 -291
rect 1181 -306 1194 -301
rect 1163 -313 1167 -310
rect 1190 -313 1194 -306
rect 1238 -313 1243 -310
rect 1065 -340 1107 -332
rect 1127 -338 1141 -331
rect 1163 -340 1167 -322
rect 1102 -356 1107 -340
rect 1164 -347 1167 -340
rect 1163 -359 1167 -347
rect 1190 -359 1194 -322
rect 1238 -342 1243 -322
rect 1211 -347 1243 -342
rect 1238 -359 1243 -347
rect 70 -369 75 -366
rect 98 -392 103 -366
rect 155 -370 160 -366
rect 357 -369 362 -366
rect -149 -404 -144 -396
rect 385 -393 390 -366
rect 442 -370 447 -366
rect 503 -368 507 -365
rect 530 -369 534 -365
rect 578 -369 583 -365
rect 702 -368 707 -365
rect 730 -395 735 -365
rect 787 -369 792 -365
rect 1017 -368 1022 -365
rect 1045 -388 1050 -365
rect 1102 -369 1107 -365
rect 1163 -367 1167 -364
rect 1190 -368 1194 -364
rect 1238 -368 1243 -364
rect -234 -431 -229 -412
rect -271 -437 -229 -431
rect -234 -452 -229 -437
rect -206 -452 -201 -412
rect -149 -428 -144 -412
rect -186 -436 -144 -428
rect -149 -452 -144 -436
rect 147 -459 152 -451
rect 175 -459 180 -451
rect 434 -459 439 -451
rect 462 -459 467 -451
rect 780 -459 785 -451
rect 808 -459 813 -451
rect 1062 -459 1067 -451
rect 1090 -459 1095 -451
rect 1389 -454 1394 -446
rect 1417 -454 1422 -446
rect -234 -464 -229 -461
rect -234 -511 -229 -503
rect -206 -511 -201 -461
rect -149 -465 -144 -461
rect 147 -484 152 -467
rect 66 -489 70 -484
rect 141 -489 152 -484
rect -149 -511 -144 -503
rect -234 -533 -229 -519
rect -262 -539 -229 -533
rect -234 -559 -229 -539
rect -206 -559 -201 -519
rect -149 -535 -144 -519
rect 66 -534 71 -489
rect 147 -507 152 -489
rect 175 -507 180 -467
rect 195 -491 200 -483
rect 434 -484 439 -467
rect 147 -519 152 -516
rect 94 -534 99 -526
rect -186 -543 -144 -535
rect -149 -559 -144 -543
rect 66 -567 71 -542
rect -234 -571 -229 -568
rect -234 -611 -229 -603
rect -206 -611 -201 -568
rect -149 -572 -144 -568
rect 47 -574 71 -567
rect 66 -582 71 -574
rect 94 -582 99 -542
rect 175 -558 180 -516
rect 233 -537 238 -491
rect 353 -489 357 -484
rect 428 -489 439 -484
rect 261 -537 266 -529
rect 353 -534 358 -489
rect 434 -507 439 -489
rect 462 -507 467 -467
rect 482 -491 487 -483
rect 780 -484 785 -467
rect 434 -519 439 -516
rect 381 -534 386 -526
rect 114 -566 180 -558
rect 66 -594 71 -591
rect -149 -611 -144 -603
rect -234 -633 -229 -619
rect -253 -639 -229 -633
rect -234 -659 -229 -639
rect -206 -659 -201 -619
rect -149 -635 -144 -619
rect -186 -643 -144 -635
rect -149 -659 -144 -643
rect 94 -639 99 -591
rect 147 -619 152 -611
rect 175 -619 180 -566
rect 233 -585 238 -545
rect 261 -585 266 -545
rect 281 -567 334 -561
rect 353 -567 358 -542
rect 281 -569 326 -567
rect 334 -574 358 -567
rect 353 -582 358 -574
rect 381 -582 386 -542
rect 462 -558 467 -516
rect 520 -537 525 -491
rect 699 -489 703 -484
rect 774 -489 785 -484
rect 548 -537 553 -529
rect 699 -534 704 -489
rect 780 -507 785 -489
rect 808 -507 813 -467
rect 828 -491 833 -483
rect 1062 -484 1067 -467
rect 780 -519 785 -516
rect 727 -534 732 -526
rect 401 -566 467 -558
rect 353 -594 358 -591
rect 233 -597 238 -594
rect 94 -656 98 -639
rect 94 -660 115 -656
rect -234 -671 -229 -668
rect -206 -671 -201 -668
rect -149 -672 -144 -668
rect 111 -712 115 -660
rect 147 -667 152 -627
rect 175 -667 180 -627
rect 261 -643 266 -594
rect 195 -651 266 -643
rect 381 -639 386 -591
rect 434 -619 439 -611
rect 462 -619 467 -566
rect 520 -585 525 -545
rect 548 -585 553 -545
rect 568 -569 619 -561
rect 699 -567 704 -542
rect 680 -574 704 -567
rect 699 -582 704 -574
rect 727 -582 732 -542
rect 808 -558 813 -516
rect 866 -537 871 -491
rect 981 -489 985 -484
rect 1056 -489 1067 -484
rect 894 -537 899 -529
rect 981 -534 986 -489
rect 1062 -507 1067 -489
rect 1090 -507 1095 -467
rect 1389 -479 1394 -462
rect 1110 -491 1115 -483
rect 1062 -519 1067 -516
rect 1009 -534 1014 -526
rect 747 -566 813 -558
rect 699 -594 704 -591
rect 520 -597 525 -594
rect 381 -656 385 -639
rect 381 -660 402 -656
rect 147 -679 152 -676
rect 175 -679 180 -676
rect 398 -712 402 -660
rect 434 -667 439 -627
rect 462 -667 467 -627
rect 548 -643 553 -594
rect 482 -651 553 -643
rect 727 -639 732 -591
rect 780 -619 785 -611
rect 808 -619 813 -566
rect 866 -585 871 -545
rect 894 -585 899 -545
rect 914 -567 962 -561
rect 981 -567 986 -542
rect 914 -569 954 -567
rect 962 -574 986 -567
rect 981 -582 986 -574
rect 1009 -582 1014 -542
rect 1090 -558 1095 -516
rect 1148 -537 1153 -491
rect 1308 -484 1312 -479
rect 1383 -484 1394 -479
rect 1308 -529 1313 -484
rect 1389 -502 1394 -484
rect 1417 -502 1422 -462
rect 1437 -486 1442 -478
rect 1389 -514 1394 -511
rect 1336 -529 1341 -521
rect 1176 -537 1181 -529
rect 1029 -566 1095 -558
rect 981 -594 986 -591
rect 866 -597 871 -594
rect 727 -656 731 -639
rect 727 -660 748 -656
rect 434 -679 439 -676
rect 462 -679 467 -676
rect 477 -708 527 -701
rect 98 -717 115 -712
rect 385 -717 402 -712
rect -235 -726 -230 -718
rect -207 -726 -202 -718
rect -150 -726 -145 -718
rect 70 -725 75 -717
rect 98 -725 103 -717
rect 155 -725 160 -717
rect 357 -725 362 -717
rect 385 -725 390 -717
rect 442 -725 447 -717
rect -235 -747 -230 -734
rect -280 -753 -230 -747
rect -235 -774 -230 -753
rect -207 -774 -202 -734
rect -150 -750 -145 -734
rect -187 -758 -145 -750
rect 70 -756 75 -733
rect -150 -774 -145 -758
rect 47 -763 75 -756
rect 70 -773 75 -763
rect 98 -773 103 -733
rect 155 -749 160 -733
rect 118 -757 160 -749
rect 357 -756 362 -733
rect 155 -773 160 -757
rect 334 -763 362 -756
rect 357 -773 362 -763
rect 385 -773 390 -733
rect 442 -749 447 -733
rect 477 -748 482 -708
rect 521 -718 527 -708
rect 744 -712 748 -660
rect 780 -667 785 -627
rect 808 -667 813 -627
rect 894 -643 899 -594
rect 828 -651 899 -643
rect 1009 -639 1014 -591
rect 1062 -619 1067 -611
rect 1090 -619 1095 -566
rect 1148 -585 1153 -545
rect 1176 -585 1181 -545
rect 1308 -561 1313 -537
rect 1196 -569 1246 -561
rect 1289 -569 1313 -561
rect 1308 -577 1313 -569
rect 1336 -577 1341 -537
rect 1417 -553 1422 -511
rect 1475 -532 1480 -486
rect 1503 -532 1508 -524
rect 1356 -561 1422 -553
rect 1308 -589 1313 -586
rect 1148 -597 1153 -594
rect 1009 -656 1013 -639
rect 1009 -660 1030 -656
rect 780 -679 785 -676
rect 808 -679 813 -676
rect 1026 -712 1030 -660
rect 1062 -667 1067 -627
rect 1090 -667 1095 -627
rect 1176 -643 1181 -594
rect 1110 -651 1181 -643
rect 1336 -634 1341 -586
rect 1389 -614 1394 -606
rect 1417 -614 1422 -561
rect 1475 -580 1480 -540
rect 1503 -580 1508 -540
rect 1523 -564 1531 -556
rect 1475 -592 1480 -589
rect 1336 -651 1340 -634
rect 1336 -655 1357 -651
rect 1062 -679 1067 -676
rect 1090 -679 1095 -676
rect 1104 -707 1155 -700
rect 1353 -707 1357 -655
rect 1389 -662 1394 -622
rect 1417 -662 1422 -622
rect 1503 -638 1508 -589
rect 1437 -646 1508 -638
rect 1389 -674 1394 -671
rect 1417 -674 1422 -671
rect 731 -717 748 -712
rect 1013 -717 1030 -712
rect 521 -723 534 -718
rect 503 -730 507 -727
rect 530 -730 534 -723
rect 703 -725 708 -717
rect 731 -725 736 -717
rect 788 -725 793 -717
rect 985 -725 990 -717
rect 1013 -725 1018 -717
rect 1070 -725 1075 -717
rect 578 -730 583 -727
rect 405 -757 447 -749
rect 467 -755 482 -748
rect 503 -757 507 -739
rect 442 -773 447 -757
rect 504 -764 507 -757
rect 503 -776 507 -764
rect 530 -776 534 -739
rect 578 -759 583 -739
rect 703 -756 708 -733
rect 551 -764 583 -759
rect 680 -763 708 -756
rect 578 -776 583 -764
rect 703 -773 708 -763
rect 731 -773 736 -733
rect 788 -749 793 -733
rect 751 -757 793 -749
rect 985 -756 990 -733
rect 788 -773 793 -757
rect 962 -763 990 -756
rect 985 -773 990 -763
rect 1013 -773 1018 -733
rect 1070 -749 1075 -733
rect 1104 -748 1109 -707
rect 1149 -718 1155 -707
rect 1340 -712 1357 -707
rect 1149 -723 1162 -718
rect 1312 -720 1317 -712
rect 1340 -720 1345 -712
rect 1397 -720 1402 -712
rect 1131 -730 1135 -727
rect 1158 -730 1162 -723
rect 1206 -730 1211 -727
rect 1033 -757 1075 -749
rect 1095 -755 1109 -748
rect 1131 -757 1135 -739
rect 1070 -773 1075 -757
rect 1132 -764 1135 -757
rect -235 -786 -230 -783
rect -235 -826 -230 -818
rect -207 -826 -202 -783
rect -150 -787 -145 -783
rect 70 -785 75 -782
rect 98 -812 103 -782
rect 155 -786 160 -782
rect 357 -785 362 -782
rect -150 -826 -145 -818
rect 385 -814 390 -782
rect 442 -786 447 -782
rect 503 -784 507 -781
rect 530 -785 534 -781
rect 578 -785 583 -781
rect 1131 -776 1135 -764
rect 1158 -776 1162 -739
rect 1206 -759 1211 -739
rect 1312 -751 1317 -728
rect 1289 -758 1317 -751
rect 1179 -764 1211 -759
rect 1206 -776 1211 -764
rect 1312 -768 1317 -758
rect 1340 -768 1345 -728
rect 1397 -744 1402 -728
rect 1360 -752 1402 -744
rect 1397 -768 1402 -752
rect 1312 -780 1317 -777
rect 703 -785 708 -782
rect 731 -812 736 -782
rect 788 -786 793 -782
rect 985 -785 990 -782
rect 1013 -812 1018 -782
rect 1070 -786 1075 -782
rect 1131 -784 1135 -781
rect 1158 -785 1162 -781
rect 1206 -785 1211 -781
rect 1340 -799 1345 -777
rect 1397 -781 1402 -777
rect -235 -850 -230 -834
rect -271 -856 -230 -850
rect -235 -874 -230 -856
rect -207 -874 -202 -834
rect -150 -850 -145 -834
rect -187 -858 -145 -850
rect -150 -874 -145 -858
rect -235 -886 -230 -883
rect -235 -933 -230 -925
rect -207 -933 -202 -883
rect -150 -887 -145 -883
rect 147 -917 152 -909
rect 175 -917 180 -909
rect 446 -917 451 -909
rect 474 -917 479 -909
rect 761 -917 766 -909
rect 789 -917 794 -909
rect 1090 -911 1095 -903
rect 1118 -911 1123 -903
rect 1405 -911 1410 -903
rect 1433 -911 1438 -903
rect -150 -933 -145 -925
rect -235 -952 -230 -941
rect -262 -958 -230 -952
rect -235 -981 -230 -958
rect -207 -981 -202 -941
rect -150 -957 -145 -941
rect -187 -965 -145 -957
rect -150 -981 -145 -965
rect -235 -993 -230 -990
rect -235 -1033 -230 -1025
rect -207 -1033 -202 -990
rect -150 -994 -145 -990
rect 66 -992 71 -947
rect 94 -992 99 -937
rect 147 -942 152 -925
rect 141 -947 152 -942
rect 147 -965 152 -947
rect 175 -965 180 -925
rect 195 -949 200 -941
rect 446 -942 451 -925
rect 147 -977 152 -974
rect 66 -1025 71 -1000
rect -150 -1033 -145 -1025
rect 47 -1032 71 -1025
rect 66 -1040 71 -1032
rect 94 -1040 99 -1000
rect 175 -1016 180 -974
rect 233 -995 238 -949
rect 440 -947 451 -942
rect 261 -995 266 -987
rect 365 -992 370 -947
rect 446 -965 451 -947
rect 474 -965 479 -925
rect 494 -949 499 -941
rect 761 -942 766 -925
rect 446 -977 451 -974
rect 393 -992 398 -984
rect 114 -1024 180 -1016
rect -235 -1052 -230 -1041
rect -253 -1058 -230 -1052
rect -235 -1081 -230 -1058
rect -207 -1081 -202 -1041
rect -150 -1057 -145 -1041
rect 66 -1052 71 -1049
rect -187 -1065 -145 -1057
rect -150 -1081 -145 -1065
rect -235 -1093 -230 -1090
rect -207 -1093 -202 -1090
rect -150 -1094 -145 -1090
rect 94 -1097 99 -1049
rect 147 -1077 152 -1069
rect 175 -1077 180 -1024
rect 233 -1043 238 -1003
rect 261 -1043 266 -1003
rect 365 -1019 370 -1000
rect 281 -1027 338 -1019
rect 346 -1027 370 -1019
rect 365 -1040 370 -1027
rect 393 -1040 398 -1000
rect 474 -1016 479 -974
rect 532 -995 537 -949
rect 680 -947 684 -942
rect 755 -947 766 -942
rect 560 -995 565 -987
rect 680 -992 685 -947
rect 761 -965 766 -947
rect 789 -965 794 -925
rect 1090 -936 1095 -919
rect 1009 -941 1013 -936
rect 1084 -941 1095 -936
rect 809 -949 814 -941
rect 761 -977 766 -974
rect 708 -992 713 -984
rect 413 -1024 479 -1016
rect 365 -1052 370 -1049
rect 233 -1055 238 -1052
rect 94 -1114 98 -1097
rect 94 -1118 115 -1114
rect -235 -1136 -230 -1128
rect -207 -1136 -202 -1128
rect -150 -1136 -145 -1128
rect -235 -1159 -230 -1144
rect -280 -1165 -230 -1159
rect -235 -1184 -230 -1165
rect -207 -1184 -202 -1144
rect -150 -1160 -145 -1144
rect -187 -1168 -145 -1160
rect -150 -1184 -145 -1168
rect 111 -1170 115 -1118
rect 147 -1125 152 -1085
rect 175 -1125 180 -1085
rect 261 -1101 266 -1052
rect 195 -1109 266 -1101
rect 393 -1097 398 -1049
rect 446 -1077 451 -1069
rect 474 -1077 479 -1024
rect 532 -1043 537 -1003
rect 560 -1043 565 -1003
rect 580 -1025 661 -1019
rect 680 -1025 685 -1000
rect 580 -1027 653 -1025
rect 661 -1032 685 -1025
rect 680 -1040 685 -1032
rect 708 -1040 713 -1000
rect 789 -1016 794 -974
rect 847 -995 852 -949
rect 1009 -986 1014 -941
rect 1090 -959 1095 -941
rect 1118 -959 1123 -919
rect 1138 -943 1143 -935
rect 1405 -936 1410 -919
rect 1090 -971 1095 -968
rect 1037 -986 1042 -978
rect 875 -995 880 -987
rect 728 -1024 794 -1016
rect 680 -1052 685 -1049
rect 532 -1055 537 -1052
rect 393 -1114 397 -1097
rect 393 -1118 414 -1114
rect 147 -1137 152 -1134
rect 175 -1137 180 -1134
rect 410 -1170 414 -1118
rect 446 -1125 451 -1085
rect 474 -1125 479 -1085
rect 560 -1101 565 -1052
rect 494 -1109 565 -1101
rect 708 -1097 713 -1049
rect 761 -1077 766 -1069
rect 789 -1077 794 -1024
rect 847 -1043 852 -1003
rect 875 -1043 880 -1003
rect 1009 -1019 1014 -994
rect 895 -1027 954 -1019
rect 990 -1026 1014 -1019
rect 1009 -1034 1014 -1026
rect 1037 -1034 1042 -994
rect 1118 -1010 1123 -968
rect 1176 -989 1181 -943
rect 1324 -941 1328 -936
rect 1399 -941 1410 -936
rect 1204 -989 1209 -981
rect 1324 -986 1329 -941
rect 1405 -959 1410 -941
rect 1433 -959 1438 -919
rect 1405 -971 1410 -968
rect 1352 -986 1357 -978
rect 1057 -1018 1123 -1010
rect 1009 -1046 1014 -1043
rect 847 -1055 852 -1052
rect 708 -1114 712 -1097
rect 708 -1118 729 -1114
rect 446 -1137 451 -1134
rect 474 -1137 479 -1134
rect 725 -1170 729 -1118
rect 761 -1125 766 -1085
rect 789 -1125 794 -1085
rect 875 -1101 880 -1052
rect 809 -1109 880 -1101
rect 1037 -1091 1042 -1043
rect 1090 -1071 1095 -1063
rect 1118 -1071 1123 -1018
rect 1176 -1037 1181 -997
rect 1204 -1037 1209 -997
rect 1224 -1019 1305 -1013
rect 1324 -1019 1329 -994
rect 1224 -1021 1297 -1019
rect 1305 -1026 1329 -1019
rect 1324 -1034 1329 -1026
rect 1352 -1034 1357 -994
rect 1433 -1010 1438 -968
rect 1491 -989 1496 -943
rect 1519 -989 1524 -981
rect 1372 -1018 1438 -1010
rect 1324 -1046 1329 -1043
rect 1176 -1049 1181 -1046
rect 1037 -1108 1041 -1091
rect 1037 -1112 1058 -1108
rect 761 -1137 766 -1134
rect 789 -1137 794 -1134
rect 1054 -1164 1058 -1112
rect 1090 -1119 1095 -1079
rect 1118 -1119 1123 -1079
rect 1204 -1095 1209 -1046
rect 1138 -1103 1209 -1095
rect 1352 -1091 1357 -1043
rect 1405 -1071 1410 -1063
rect 1433 -1071 1438 -1018
rect 1491 -1037 1496 -997
rect 1519 -1037 1524 -997
rect 1539 -1021 1547 -1013
rect 1491 -1049 1496 -1046
rect 1352 -1108 1356 -1091
rect 1352 -1112 1373 -1108
rect 1090 -1131 1095 -1128
rect 1118 -1131 1123 -1128
rect 1369 -1164 1373 -1112
rect 1405 -1119 1410 -1079
rect 1433 -1119 1438 -1079
rect 1519 -1095 1524 -1046
rect 1453 -1103 1524 -1095
rect 1405 -1131 1410 -1128
rect 1433 -1131 1438 -1128
rect 1041 -1169 1058 -1164
rect 1356 -1169 1373 -1164
rect 98 -1175 115 -1170
rect 397 -1175 414 -1170
rect 712 -1175 729 -1170
rect 70 -1183 75 -1175
rect 98 -1183 103 -1175
rect 155 -1183 160 -1175
rect 369 -1183 374 -1175
rect 397 -1183 402 -1175
rect 454 -1183 459 -1175
rect 684 -1183 689 -1175
rect 712 -1183 717 -1175
rect 769 -1183 774 -1175
rect 804 -1178 854 -1171
rect 1013 -1177 1018 -1169
rect 1041 -1177 1046 -1169
rect 1098 -1177 1103 -1169
rect 1328 -1177 1333 -1169
rect 1356 -1177 1361 -1169
rect 1413 -1177 1418 -1169
rect 1448 -1172 1498 -1165
rect -235 -1196 -230 -1193
rect -235 -1236 -230 -1228
rect -207 -1236 -202 -1193
rect -150 -1197 -145 -1193
rect 70 -1214 75 -1191
rect 47 -1221 75 -1214
rect -150 -1236 -145 -1228
rect 70 -1231 75 -1221
rect 98 -1231 103 -1191
rect 155 -1207 160 -1191
rect 118 -1215 160 -1207
rect 369 -1214 374 -1191
rect 155 -1231 160 -1215
rect 346 -1221 374 -1214
rect 369 -1231 374 -1221
rect 397 -1231 402 -1191
rect 454 -1207 459 -1191
rect 417 -1215 459 -1207
rect 684 -1214 689 -1191
rect 454 -1231 459 -1215
rect 661 -1221 689 -1214
rect 684 -1231 689 -1221
rect 712 -1231 717 -1191
rect 769 -1207 774 -1191
rect 804 -1206 809 -1178
rect 848 -1196 854 -1178
rect 848 -1201 861 -1196
rect 732 -1215 774 -1207
rect 794 -1213 809 -1206
rect 830 -1208 834 -1205
rect 857 -1208 861 -1201
rect 905 -1208 910 -1205
rect 1013 -1208 1018 -1185
rect 769 -1231 774 -1215
rect 990 -1215 1018 -1208
rect 830 -1235 834 -1217
rect 70 -1243 75 -1240
rect 98 -1243 103 -1240
rect 155 -1244 160 -1240
rect 369 -1243 374 -1240
rect -235 -1262 -230 -1244
rect -271 -1268 -230 -1262
rect -235 -1284 -230 -1268
rect -207 -1284 -202 -1244
rect -150 -1260 -145 -1244
rect -187 -1268 -145 -1260
rect 397 -1260 402 -1240
rect 454 -1244 459 -1240
rect 684 -1243 689 -1240
rect -150 -1284 -145 -1268
rect 712 -1278 717 -1240
rect 769 -1244 774 -1240
rect 831 -1242 834 -1235
rect 830 -1254 834 -1242
rect 857 -1254 861 -1217
rect 905 -1237 910 -1217
rect 1013 -1225 1018 -1215
rect 1041 -1225 1046 -1185
rect 1098 -1201 1103 -1185
rect 1061 -1209 1103 -1201
rect 1328 -1208 1333 -1185
rect 1098 -1225 1103 -1209
rect 1305 -1215 1333 -1208
rect 1328 -1225 1333 -1215
rect 1356 -1225 1361 -1185
rect 1413 -1201 1418 -1185
rect 1448 -1200 1453 -1172
rect 1492 -1190 1498 -1172
rect 1492 -1195 1505 -1190
rect 1376 -1209 1418 -1201
rect 1438 -1207 1453 -1200
rect 1474 -1202 1478 -1199
rect 1501 -1202 1505 -1195
rect 1549 -1202 1554 -1199
rect 1413 -1225 1418 -1209
rect 1474 -1229 1478 -1211
rect 1013 -1237 1018 -1234
rect 878 -1242 910 -1237
rect 905 -1254 910 -1242
rect 830 -1262 834 -1259
rect 857 -1263 861 -1259
rect 905 -1263 910 -1259
rect 1041 -1264 1046 -1234
rect 1098 -1238 1103 -1234
rect 1328 -1237 1333 -1234
rect 1356 -1274 1361 -1234
rect 1413 -1238 1418 -1234
rect 1475 -1236 1478 -1229
rect 1474 -1248 1478 -1236
rect 1501 -1248 1505 -1211
rect 1549 -1231 1554 -1211
rect 1522 -1236 1554 -1231
rect 1549 -1248 1554 -1236
rect 1474 -1256 1478 -1253
rect 1501 -1257 1505 -1253
rect 1549 -1257 1554 -1253
rect 147 -1291 152 -1283
rect 175 -1291 180 -1283
rect -235 -1296 -230 -1293
rect -235 -1343 -230 -1335
rect -207 -1343 -202 -1293
rect -150 -1297 -145 -1293
rect 66 -1321 70 -1316
rect -150 -1343 -145 -1335
rect -235 -1364 -230 -1351
rect -262 -1370 -230 -1364
rect -235 -1391 -230 -1370
rect -207 -1391 -202 -1351
rect -150 -1367 -145 -1351
rect 66 -1366 71 -1321
rect 94 -1366 99 -1313
rect 147 -1316 152 -1299
rect 141 -1321 152 -1316
rect 147 -1339 152 -1321
rect 175 -1339 180 -1299
rect 195 -1323 200 -1315
rect 147 -1351 152 -1348
rect -187 -1375 -145 -1367
rect -150 -1391 -145 -1375
rect 66 -1399 71 -1374
rect -235 -1403 -230 -1400
rect -235 -1443 -230 -1435
rect -207 -1443 -202 -1400
rect -150 -1404 -145 -1400
rect 47 -1406 71 -1399
rect 66 -1414 71 -1406
rect 94 -1414 99 -1374
rect 175 -1390 180 -1348
rect 233 -1369 238 -1323
rect 478 -1324 483 -1316
rect 506 -1324 511 -1316
rect 793 -1324 798 -1316
rect 821 -1324 826 -1316
rect 478 -1349 483 -1332
rect 397 -1354 401 -1349
rect 472 -1354 483 -1349
rect 261 -1369 266 -1361
rect 114 -1398 180 -1390
rect 66 -1426 71 -1423
rect -150 -1443 -145 -1435
rect -235 -1464 -230 -1451
rect -253 -1470 -230 -1464
rect -235 -1491 -230 -1470
rect -207 -1491 -202 -1451
rect -150 -1467 -145 -1451
rect -187 -1475 -145 -1467
rect -150 -1491 -145 -1475
rect 94 -1471 99 -1423
rect 147 -1451 152 -1443
rect 175 -1451 180 -1398
rect 233 -1417 238 -1377
rect 261 -1417 266 -1377
rect 397 -1399 402 -1354
rect 478 -1372 483 -1354
rect 506 -1372 511 -1332
rect 526 -1356 531 -1348
rect 793 -1349 798 -1332
rect 478 -1384 483 -1381
rect 425 -1399 430 -1391
rect 233 -1429 238 -1426
rect 94 -1488 98 -1471
rect 94 -1492 115 -1488
rect -235 -1503 -230 -1500
rect -207 -1503 -202 -1500
rect -150 -1504 -145 -1500
rect 111 -1544 115 -1492
rect 147 -1499 152 -1459
rect 175 -1499 180 -1459
rect 261 -1475 266 -1426
rect 397 -1432 402 -1407
rect 378 -1439 402 -1432
rect 397 -1447 402 -1439
rect 425 -1447 430 -1407
rect 506 -1423 511 -1381
rect 564 -1402 569 -1356
rect 712 -1354 716 -1349
rect 787 -1354 798 -1349
rect 592 -1402 597 -1394
rect 712 -1399 717 -1354
rect 793 -1372 798 -1354
rect 821 -1372 826 -1332
rect 841 -1356 846 -1348
rect 793 -1384 798 -1381
rect 740 -1399 745 -1391
rect 445 -1431 511 -1423
rect 397 -1459 402 -1456
rect 195 -1483 266 -1475
rect 425 -1504 430 -1456
rect 478 -1484 483 -1476
rect 506 -1484 511 -1431
rect 564 -1450 569 -1410
rect 592 -1450 597 -1410
rect 612 -1432 693 -1426
rect 712 -1432 717 -1407
rect 612 -1434 685 -1432
rect 693 -1439 717 -1432
rect 712 -1447 717 -1439
rect 740 -1447 745 -1407
rect 821 -1423 826 -1381
rect 879 -1402 884 -1356
rect 907 -1402 912 -1394
rect 760 -1431 826 -1423
rect 712 -1459 717 -1456
rect 564 -1462 569 -1459
rect 147 -1511 152 -1508
rect 175 -1511 180 -1508
rect 425 -1521 429 -1504
rect 425 -1525 446 -1521
rect 98 -1549 115 -1544
rect 70 -1557 75 -1549
rect 98 -1557 103 -1549
rect 155 -1557 160 -1549
rect 70 -1588 75 -1565
rect 47 -1595 75 -1588
rect 70 -1605 75 -1595
rect 98 -1605 103 -1565
rect 155 -1581 160 -1565
rect 442 -1577 446 -1525
rect 478 -1532 483 -1492
rect 506 -1532 511 -1492
rect 592 -1508 597 -1459
rect 526 -1516 597 -1508
rect 740 -1504 745 -1456
rect 793 -1484 798 -1476
rect 821 -1484 826 -1431
rect 879 -1450 884 -1410
rect 907 -1450 912 -1410
rect 927 -1434 935 -1426
rect 879 -1462 884 -1459
rect 740 -1521 744 -1504
rect 740 -1525 761 -1521
rect 478 -1544 483 -1541
rect 506 -1544 511 -1541
rect 757 -1577 761 -1525
rect 793 -1532 798 -1492
rect 821 -1532 826 -1492
rect 907 -1508 912 -1459
rect 841 -1516 912 -1508
rect 793 -1544 798 -1541
rect 821 -1544 826 -1541
rect 118 -1589 160 -1581
rect 429 -1582 446 -1577
rect 744 -1582 761 -1577
rect 155 -1605 160 -1589
rect 401 -1590 406 -1582
rect 429 -1590 434 -1582
rect 486 -1590 491 -1582
rect 716 -1590 721 -1582
rect 744 -1590 749 -1582
rect 801 -1590 806 -1582
rect 836 -1585 886 -1578
rect 70 -1617 75 -1614
rect 98 -1617 103 -1614
rect 155 -1618 160 -1614
rect 401 -1621 406 -1598
rect 378 -1628 406 -1621
rect 401 -1638 406 -1628
rect 429 -1638 434 -1598
rect 486 -1614 491 -1598
rect 449 -1622 491 -1614
rect 716 -1621 721 -1598
rect 486 -1638 491 -1622
rect 693 -1628 721 -1621
rect 716 -1638 721 -1628
rect 744 -1638 749 -1598
rect 801 -1614 806 -1598
rect 836 -1613 841 -1585
rect 880 -1603 886 -1585
rect 880 -1608 893 -1603
rect 764 -1622 806 -1614
rect 826 -1620 841 -1613
rect 862 -1615 866 -1612
rect 889 -1615 893 -1608
rect 937 -1615 942 -1612
rect 801 -1638 806 -1622
rect 862 -1642 866 -1624
rect 401 -1650 406 -1647
rect 147 -1667 152 -1659
rect 175 -1667 180 -1659
rect 66 -1697 70 -1692
rect 66 -1742 71 -1697
rect 94 -1742 99 -1684
rect 147 -1692 152 -1675
rect 141 -1697 152 -1692
rect 147 -1715 152 -1697
rect 175 -1715 180 -1675
rect 429 -1677 434 -1647
rect 486 -1651 491 -1647
rect 716 -1650 721 -1647
rect 744 -1686 749 -1647
rect 801 -1651 806 -1647
rect 863 -1649 866 -1642
rect 862 -1661 866 -1649
rect 889 -1661 893 -1624
rect 937 -1644 942 -1624
rect 910 -1649 942 -1644
rect 937 -1661 942 -1649
rect 862 -1669 866 -1666
rect 889 -1670 893 -1666
rect 937 -1670 942 -1666
rect 195 -1699 200 -1691
rect 147 -1727 152 -1724
rect 66 -1775 71 -1750
rect 47 -1782 71 -1775
rect 66 -1790 71 -1782
rect 94 -1790 99 -1750
rect 175 -1766 180 -1724
rect 233 -1745 238 -1699
rect 261 -1745 266 -1737
rect 114 -1774 180 -1766
rect 66 -1802 71 -1799
rect 94 -1847 99 -1799
rect 147 -1827 152 -1819
rect 175 -1827 180 -1774
rect 233 -1793 238 -1753
rect 261 -1793 266 -1753
rect 281 -1777 289 -1769
rect 233 -1805 238 -1802
rect 94 -1864 98 -1847
rect 94 -1868 115 -1864
rect 111 -1920 115 -1868
rect 147 -1875 152 -1835
rect 175 -1875 180 -1835
rect 261 -1851 266 -1802
rect 195 -1859 266 -1851
rect 147 -1887 152 -1884
rect 175 -1887 180 -1884
rect 98 -1925 115 -1920
rect 70 -1933 75 -1925
rect 98 -1933 103 -1925
rect 155 -1933 160 -1925
rect 70 -1964 75 -1941
rect 47 -1971 75 -1964
rect 70 -1981 75 -1971
rect 98 -1981 103 -1941
rect 155 -1957 160 -1941
rect 118 -1965 160 -1957
rect 155 -1981 160 -1965
rect 70 -1993 75 -1990
rect 98 -1993 103 -1990
rect 155 -1994 160 -1990
<< polycontact >>
rect 70 330 74 335
rect 137 330 141 335
rect 381 343 386 350
rect 187 328 195 336
rect 200 328 207 336
rect 232 328 238 336
rect 39 245 47 252
rect 357 330 361 335
rect 424 330 428 335
rect 474 328 482 336
rect 487 328 494 336
rect 519 328 525 336
rect 106 253 114 261
rect 273 250 281 258
rect 326 245 334 252
rect 393 253 401 261
rect 98 174 103 180
rect 142 174 147 180
rect 187 168 195 176
rect 560 250 568 258
rect 385 174 390 180
rect 429 174 434 180
rect 474 168 482 176
rect -286 68 -280 74
rect -194 74 -186 82
rect 39 56 47 63
rect 110 62 118 70
rect 326 56 334 63
rect 397 62 405 70
rect 462 64 467 71
rect 497 55 504 62
rect 546 55 551 60
rect 98 3 103 7
rect -277 -35 -271 -29
rect -194 -26 -186 -18
rect 70 -73 74 -68
rect 137 -73 141 -68
rect -268 -137 -262 -131
rect 187 -75 195 -67
rect 200 -75 207 -67
rect 232 -75 238 -67
rect -194 -133 -186 -125
rect 39 -158 47 -151
rect 357 -73 361 -68
rect 424 -73 428 -68
rect 474 -75 482 -67
rect 487 -75 494 -67
rect 519 -75 525 -67
rect 106 -150 114 -142
rect -259 -237 -253 -231
rect -194 -233 -186 -225
rect 273 -153 281 -145
rect 326 -158 334 -151
rect 702 -72 706 -67
rect 769 -72 773 -67
rect 819 -74 827 -66
rect 832 -74 839 -66
rect 864 -74 870 -66
rect 393 -150 401 -142
rect 98 -229 103 -223
rect 142 -229 147 -223
rect 187 -235 195 -227
rect 560 -153 568 -145
rect 619 -153 627 -145
rect 671 -157 679 -150
rect 1017 -72 1021 -67
rect 1084 -72 1088 -67
rect 1134 -74 1142 -66
rect 1147 -74 1154 -66
rect 1179 -74 1185 -66
rect 738 -149 746 -141
rect 385 -229 390 -223
rect 429 -229 434 -223
rect 474 -235 482 -227
rect 905 -152 913 -144
rect 986 -157 994 -150
rect 1053 -149 1061 -141
rect 730 -228 735 -222
rect 774 -228 779 -222
rect -286 -334 -280 -328
rect -194 -336 -186 -328
rect 39 -347 47 -340
rect 110 -341 118 -333
rect 326 -347 334 -340
rect 819 -234 827 -226
rect 1220 -152 1228 -144
rect 1045 -228 1050 -222
rect 1089 -228 1094 -222
rect 1134 -234 1142 -226
rect 397 -341 405 -333
rect 462 -339 467 -332
rect 497 -348 504 -341
rect 546 -348 551 -343
rect 671 -346 679 -339
rect 742 -340 750 -332
rect 986 -346 994 -339
rect 1057 -340 1065 -332
rect 1122 -338 1127 -331
rect 1157 -347 1164 -340
rect 1206 -347 1211 -342
rect 98 -399 103 -392
rect 385 -397 390 -393
rect 1045 -393 1050 -388
rect 730 -399 735 -395
rect -277 -437 -271 -431
rect -194 -436 -186 -428
rect 70 -489 74 -484
rect 137 -489 141 -484
rect -268 -539 -262 -533
rect 187 -491 195 -483
rect 200 -491 207 -483
rect 232 -491 238 -483
rect -194 -543 -186 -535
rect 39 -574 47 -567
rect 357 -489 361 -484
rect 424 -489 428 -484
rect 474 -491 482 -483
rect 487 -491 494 -483
rect 519 -491 525 -483
rect 106 -566 114 -558
rect -259 -639 -253 -633
rect -194 -643 -186 -635
rect 273 -569 281 -561
rect 326 -574 334 -567
rect 703 -489 707 -484
rect 770 -489 774 -484
rect 820 -491 828 -483
rect 833 -491 840 -483
rect 865 -491 871 -483
rect 393 -566 401 -558
rect 98 -645 103 -639
rect 142 -645 147 -639
rect 187 -651 195 -643
rect 560 -569 568 -561
rect 619 -569 626 -561
rect 672 -574 680 -567
rect 985 -489 989 -484
rect 1052 -489 1056 -484
rect 1102 -491 1110 -483
rect 1115 -491 1122 -483
rect 1147 -491 1153 -483
rect 739 -566 747 -558
rect 385 -645 390 -639
rect 429 -645 434 -639
rect 474 -651 482 -643
rect 906 -569 914 -561
rect 954 -574 962 -567
rect 1312 -484 1316 -479
rect 1379 -484 1383 -479
rect 1429 -486 1437 -478
rect 1442 -486 1449 -478
rect 1474 -486 1480 -478
rect 1021 -566 1029 -558
rect 731 -645 736 -639
rect 775 -645 780 -639
rect -286 -753 -280 -747
rect -195 -758 -187 -750
rect 39 -763 47 -756
rect 110 -757 118 -749
rect 326 -763 334 -756
rect 820 -651 828 -643
rect 1188 -569 1196 -561
rect 1246 -569 1253 -561
rect 1281 -569 1289 -561
rect 1348 -561 1356 -553
rect 1013 -645 1018 -639
rect 1057 -645 1062 -639
rect 1102 -651 1110 -643
rect 1515 -564 1523 -556
rect 1340 -640 1345 -634
rect 1384 -640 1389 -634
rect 1429 -646 1437 -638
rect 397 -757 405 -749
rect 462 -755 467 -748
rect 497 -764 504 -757
rect 546 -764 551 -759
rect 672 -763 680 -756
rect 743 -757 751 -749
rect 954 -763 962 -756
rect 1025 -757 1033 -749
rect 1090 -755 1095 -748
rect 1125 -764 1132 -757
rect 98 -819 103 -812
rect 1281 -758 1289 -751
rect 1174 -764 1179 -759
rect 1352 -752 1360 -744
rect 385 -822 390 -814
rect 731 -816 736 -812
rect 1340 -806 1345 -799
rect 1013 -820 1018 -812
rect -277 -856 -271 -850
rect -195 -858 -187 -850
rect 94 -937 99 -930
rect -268 -958 -262 -952
rect -195 -965 -187 -957
rect 66 -947 71 -942
rect 137 -947 141 -942
rect 187 -949 195 -941
rect 200 -949 207 -941
rect 232 -949 238 -941
rect 39 -1032 47 -1025
rect 365 -947 370 -942
rect 436 -947 440 -942
rect 486 -949 494 -941
rect 499 -949 506 -941
rect 531 -949 537 -941
rect 106 -1024 114 -1016
rect -259 -1058 -253 -1052
rect -195 -1065 -187 -1057
rect 273 -1027 281 -1019
rect 338 -1027 346 -1019
rect 684 -947 688 -942
rect 751 -947 755 -942
rect 1013 -941 1017 -936
rect 1080 -941 1084 -936
rect 801 -949 809 -941
rect 814 -949 821 -941
rect 846 -949 852 -941
rect 405 -1024 413 -1016
rect 98 -1103 103 -1097
rect 142 -1103 147 -1097
rect -286 -1165 -280 -1159
rect -195 -1168 -187 -1160
rect 187 -1109 195 -1101
rect 572 -1027 580 -1019
rect 653 -1032 661 -1025
rect 1130 -943 1138 -935
rect 1143 -943 1150 -935
rect 1175 -943 1181 -935
rect 720 -1024 728 -1016
rect 397 -1103 402 -1097
rect 441 -1103 446 -1097
rect 486 -1109 494 -1101
rect 887 -1027 895 -1019
rect 954 -1027 962 -1019
rect 982 -1026 990 -1019
rect 1328 -941 1332 -936
rect 1395 -941 1399 -936
rect 1490 -943 1496 -935
rect 1049 -1018 1057 -1010
rect 712 -1103 717 -1097
rect 756 -1103 761 -1097
rect 801 -1109 809 -1101
rect 1216 -1021 1224 -1013
rect 1297 -1026 1305 -1019
rect 1364 -1018 1372 -1010
rect 1041 -1097 1046 -1091
rect 1085 -1097 1090 -1091
rect 1130 -1103 1138 -1095
rect 1531 -1021 1539 -1013
rect 1356 -1097 1361 -1091
rect 1400 -1097 1405 -1091
rect 1445 -1103 1453 -1095
rect 39 -1221 47 -1214
rect 110 -1215 118 -1207
rect 338 -1221 346 -1214
rect 409 -1215 417 -1207
rect 653 -1221 661 -1214
rect 724 -1215 732 -1207
rect 789 -1213 794 -1206
rect 982 -1215 990 -1208
rect -277 -1268 -271 -1262
rect -195 -1268 -187 -1260
rect 397 -1266 402 -1260
rect 824 -1242 831 -1235
rect 1053 -1209 1061 -1201
rect 1297 -1215 1305 -1208
rect 1368 -1209 1376 -1201
rect 1433 -1207 1438 -1200
rect 873 -1242 878 -1237
rect 1041 -1268 1046 -1264
rect 1468 -1236 1475 -1229
rect 1517 -1236 1522 -1231
rect 712 -1286 717 -1278
rect 1356 -1279 1361 -1274
rect 94 -1313 99 -1307
rect 70 -1321 74 -1316
rect -268 -1370 -262 -1364
rect 137 -1321 141 -1316
rect 187 -1323 195 -1315
rect 200 -1323 207 -1315
rect 232 -1323 238 -1315
rect -195 -1375 -187 -1367
rect 39 -1406 47 -1399
rect 401 -1354 405 -1349
rect 468 -1354 472 -1349
rect 106 -1398 114 -1390
rect -259 -1470 -253 -1464
rect -195 -1475 -187 -1467
rect 273 -1401 281 -1393
rect 518 -1356 526 -1348
rect 531 -1356 538 -1348
rect 563 -1356 569 -1348
rect 98 -1477 103 -1471
rect 142 -1477 147 -1471
rect 370 -1439 378 -1432
rect 716 -1354 720 -1349
rect 783 -1354 787 -1349
rect 833 -1356 841 -1348
rect 846 -1356 853 -1348
rect 878 -1356 884 -1348
rect 437 -1431 445 -1423
rect 187 -1483 195 -1475
rect 604 -1434 612 -1426
rect 685 -1439 693 -1432
rect 752 -1431 760 -1423
rect 429 -1510 434 -1504
rect 473 -1510 478 -1504
rect 39 -1595 47 -1588
rect 518 -1516 526 -1508
rect 919 -1434 927 -1426
rect 744 -1510 749 -1504
rect 788 -1510 793 -1504
rect 833 -1516 841 -1508
rect 110 -1589 118 -1581
rect 370 -1628 378 -1621
rect 441 -1622 449 -1614
rect 685 -1628 693 -1621
rect 756 -1622 764 -1614
rect 821 -1620 826 -1613
rect 94 -1684 99 -1679
rect 70 -1697 74 -1692
rect 137 -1697 141 -1692
rect 429 -1684 434 -1677
rect 856 -1649 863 -1642
rect 905 -1649 910 -1644
rect 744 -1690 749 -1686
rect 187 -1699 195 -1691
rect 200 -1699 207 -1691
rect 232 -1699 238 -1691
rect 39 -1782 47 -1775
rect 106 -1774 114 -1766
rect 273 -1777 281 -1769
rect 98 -1853 103 -1847
rect 142 -1853 147 -1847
rect 187 -1859 195 -1851
rect 39 -1971 47 -1964
rect 110 -1965 118 -1957
<< metal1 >>
rect 144 375 157 382
rect 164 375 178 382
rect 185 375 197 382
rect 138 360 145 375
rect 187 360 194 375
rect 160 336 167 352
rect 381 350 386 386
rect 431 375 444 382
rect 451 375 465 382
rect 472 375 484 382
rect 425 360 432 375
rect 474 360 481 375
rect 447 336 454 352
rect 74 330 137 335
rect 160 328 187 336
rect 207 328 232 336
rect 361 330 424 335
rect 447 328 474 336
rect 494 328 519 336
rect 187 312 195 328
rect 474 312 482 328
rect 62 300 76 307
rect 83 300 97 307
rect 104 300 118 307
rect 57 285 64 300
rect 106 285 113 300
rect 133 294 141 303
rect 231 299 243 304
rect 224 297 243 299
rect 250 297 264 304
rect 271 297 289 304
rect 349 300 363 307
rect 370 300 387 307
rect 394 300 405 307
rect 133 286 145 294
rect 153 286 198 294
rect 224 282 231 297
rect 273 282 280 297
rect 79 261 86 277
rect 344 285 351 300
rect 393 285 400 300
rect 420 294 428 303
rect 518 299 530 304
rect 511 297 530 299
rect 537 297 551 304
rect 558 297 588 304
rect 420 286 432 294
rect 440 286 485 294
rect 511 282 518 297
rect 560 282 567 297
rect 79 253 106 261
rect -243 121 -224 127
rect -217 121 -200 127
rect -193 121 -151 127
rect -143 121 -133 127
rect -124 121 -119 127
rect -243 106 -236 121
rect -194 106 -187 121
rect -158 106 -151 121
rect -221 82 -214 98
rect -221 74 -194 82
rect -286 -328 -280 68
rect -194 58 -186 74
rect -136 69 -129 98
rect 39 69 47 245
rect 106 237 114 253
rect 246 258 253 274
rect 366 261 373 277
rect 246 250 273 258
rect 366 253 393 261
rect 273 234 281 250
rect 52 219 60 228
rect 58 211 64 219
rect 72 211 122 219
rect 144 215 157 222
rect 164 215 181 222
rect 188 215 203 222
rect 219 216 227 225
rect 138 200 145 215
rect 187 200 194 215
rect 228 208 231 216
rect 239 208 289 216
rect 103 174 142 180
rect 160 176 167 192
rect 160 168 187 176
rect 187 152 195 168
rect 133 135 141 143
rect 141 126 145 134
rect 153 126 173 134
rect 181 126 197 134
rect 66 109 80 115
rect 87 109 101 115
rect 108 109 153 115
rect 161 109 171 115
rect 180 109 183 115
rect 66 108 68 109
rect 61 94 68 108
rect 110 94 117 109
rect 146 94 153 109
rect -136 63 47 69
rect -136 58 -129 63
rect 83 70 90 86
rect 168 71 175 86
rect 83 62 110 70
rect -248 40 -240 49
rect -165 40 -157 49
rect 110 46 118 62
rect 168 46 175 63
rect -240 32 -236 40
rect -228 32 -200 40
rect -192 32 -157 40
rect -148 32 -138 40
rect -129 37 -128 40
rect -129 32 64 37
rect 56 28 64 32
rect 139 28 147 37
rect 186 29 195 126
rect 326 63 334 245
rect 393 237 401 253
rect 533 258 540 274
rect 533 250 560 258
rect 560 234 568 250
rect 339 219 347 228
rect 345 211 351 219
rect 359 211 409 219
rect 431 215 444 222
rect 451 215 468 222
rect 475 215 490 222
rect 506 216 514 225
rect 425 200 432 215
rect 474 200 481 215
rect 515 208 518 216
rect 526 208 576 216
rect 390 174 429 180
rect 447 176 454 192
rect 447 168 474 176
rect 474 152 482 168
rect 420 135 428 143
rect 428 126 432 134
rect 440 126 460 134
rect 468 126 484 134
rect 353 109 367 115
rect 374 109 388 115
rect 395 109 440 115
rect 448 109 458 115
rect 467 109 470 115
rect 353 108 355 109
rect 348 94 355 108
rect 397 94 404 109
rect 433 94 440 109
rect 370 70 377 86
rect 370 62 397 70
rect 397 46 405 62
rect 455 46 462 86
rect 343 29 351 37
rect 186 28 351 29
rect 426 28 434 37
rect 473 28 482 126
rect 583 110 588 297
rect 495 104 504 110
rect 510 104 530 110
rect 536 104 557 110
rect 563 104 576 110
rect 582 104 588 110
rect 495 89 500 104
rect 568 89 573 104
rect 491 55 497 62
rect 541 60 546 80
rect 514 55 546 60
rect 514 43 520 55
rect 589 43 594 80
rect -243 21 -224 27
rect -217 21 -197 27
rect -189 21 -151 27
rect -143 21 -133 27
rect -124 21 -119 27
rect -243 6 -236 21
rect -194 6 -187 21
rect -158 6 -151 21
rect 56 20 68 28
rect 76 20 105 28
rect 113 20 147 28
rect 156 20 166 28
rect 175 20 355 28
rect 363 20 383 28
rect 391 20 434 28
rect 443 20 453 28
rect 462 26 482 28
rect 494 26 499 38
rect 540 26 545 38
rect 563 26 569 38
rect 462 20 500 26
rect 506 20 531 26
rect 537 20 553 26
rect 559 20 572 26
rect 578 20 586 26
rect -221 -18 -214 -2
rect -221 -26 -194 -18
rect -286 -747 -280 -334
rect -286 -1159 -280 -753
rect -277 -431 -271 -35
rect -194 -42 -186 -26
rect -136 -20 -129 -2
rect 98 -3 103 3
rect -136 -28 -74 -20
rect 144 -28 157 -21
rect 164 -28 178 -21
rect 185 -28 197 -21
rect 431 -28 444 -21
rect 451 -28 465 -21
rect 472 -28 484 -21
rect 776 -27 789 -20
rect 796 -27 810 -20
rect 817 -27 829 -20
rect 1091 -27 1104 -20
rect 1111 -27 1125 -20
rect 1132 -27 1144 -20
rect -136 -42 -129 -28
rect 138 -43 145 -28
rect 187 -43 194 -28
rect 425 -43 432 -28
rect 474 -43 481 -28
rect 770 -42 777 -27
rect 819 -42 826 -27
rect 1085 -42 1092 -27
rect 1134 -42 1141 -27
rect -248 -60 -240 -51
rect -165 -60 -157 -51
rect -240 -68 -236 -60
rect -228 -68 -200 -60
rect -192 -68 -157 -60
rect -148 -68 -138 -60
rect -129 -68 -128 -60
rect 160 -67 167 -51
rect 447 -67 454 -51
rect 792 -66 799 -50
rect 1107 -66 1114 -50
rect 74 -73 137 -68
rect 160 -75 187 -67
rect 207 -75 232 -67
rect 361 -73 424 -68
rect 447 -75 474 -67
rect 494 -75 519 -67
rect 706 -72 769 -67
rect 792 -74 819 -66
rect 839 -74 864 -66
rect 1021 -72 1084 -67
rect 1107 -74 1134 -66
rect 1154 -74 1179 -66
rect -243 -86 -224 -80
rect -217 -86 -151 -80
rect -143 -86 -133 -80
rect -124 -86 -119 -80
rect -114 -86 62 -80
rect -243 -101 -236 -86
rect -194 -101 -187 -86
rect -158 -101 -151 -86
rect -115 -87 62 -86
rect 56 -96 62 -87
rect 187 -91 195 -75
rect 474 -91 482 -75
rect 819 -90 827 -74
rect 1134 -90 1142 -74
rect 56 -103 57 -96
rect 62 -103 76 -96
rect 83 -103 97 -96
rect 104 -103 118 -96
rect -221 -125 -214 -109
rect -277 -850 -271 -437
rect -277 -1262 -271 -856
rect -221 -133 -194 -125
rect -268 -533 -262 -137
rect -194 -149 -186 -133
rect -136 -127 -129 -109
rect 57 -118 64 -103
rect 106 -118 113 -103
rect 133 -109 141 -100
rect 231 -104 243 -99
rect 224 -106 243 -104
rect 250 -106 264 -99
rect 271 -106 289 -99
rect 349 -103 363 -96
rect 370 -103 384 -96
rect 391 -103 405 -96
rect 133 -117 145 -109
rect 153 -117 198 -109
rect 224 -121 231 -106
rect 273 -121 280 -106
rect -136 -135 -86 -127
rect -136 -149 -129 -135
rect 79 -142 86 -126
rect 344 -118 351 -103
rect 393 -118 400 -103
rect 420 -109 428 -100
rect 518 -104 530 -99
rect 511 -106 530 -104
rect 537 -106 551 -99
rect 558 -102 689 -99
rect 694 -102 708 -95
rect 715 -102 729 -95
rect 736 -102 750 -95
rect 558 -106 696 -102
rect 420 -117 432 -109
rect 440 -117 485 -109
rect 511 -121 518 -106
rect 560 -121 567 -106
rect 79 -150 106 -142
rect -248 -167 -240 -158
rect -165 -167 -157 -158
rect -240 -175 -236 -167
rect -228 -175 -200 -167
rect -192 -175 -157 -167
rect -148 -175 -138 -167
rect -129 -175 -128 -167
rect -243 -186 -224 -180
rect -217 -186 -197 -180
rect -190 -186 -151 -180
rect -143 -186 -133 -180
rect -124 -186 -119 -180
rect -243 -201 -236 -186
rect -194 -201 -187 -186
rect -158 -201 -151 -186
rect -221 -225 -214 -209
rect -268 -952 -262 -539
rect -268 -1364 -262 -958
rect -221 -233 -194 -225
rect -259 -633 -253 -237
rect -194 -249 -186 -233
rect -136 -228 -129 -209
rect -136 -235 -108 -228
rect -136 -249 -129 -235
rect -248 -267 -240 -258
rect -165 -267 -157 -258
rect -240 -275 -236 -267
rect -228 -275 -200 -267
rect -192 -275 -157 -267
rect -148 -275 -138 -267
rect -129 -275 -128 -267
rect -243 -289 -224 -283
rect -217 -289 -201 -283
rect -194 -289 -151 -283
rect -143 -289 -133 -283
rect -124 -289 -119 -283
rect -243 -304 -236 -289
rect -194 -304 -187 -289
rect -158 -304 -151 -289
rect -221 -328 -214 -312
rect -221 -336 -194 -328
rect -194 -352 -186 -336
rect -136 -331 -129 -312
rect 39 -331 47 -158
rect 106 -166 114 -150
rect 246 -145 253 -129
rect 366 -142 373 -126
rect 246 -153 273 -145
rect 366 -150 393 -142
rect 273 -169 281 -153
rect 52 -184 60 -175
rect 58 -192 64 -184
rect 72 -192 122 -184
rect 144 -188 157 -181
rect 164 -188 181 -181
rect 188 -188 203 -181
rect 219 -187 227 -178
rect 138 -203 145 -188
rect 187 -203 194 -188
rect 228 -195 231 -187
rect 239 -195 289 -187
rect 103 -229 142 -223
rect 160 -227 167 -211
rect 160 -235 187 -227
rect 187 -251 195 -235
rect 133 -268 141 -260
rect 141 -277 145 -269
rect 153 -277 173 -269
rect 181 -277 197 -269
rect 66 -294 80 -288
rect 87 -294 101 -288
rect 108 -294 153 -288
rect 161 -294 171 -288
rect 180 -294 183 -288
rect 66 -295 68 -294
rect 61 -309 68 -295
rect 110 -309 117 -294
rect 146 -309 153 -294
rect -136 -338 47 -331
rect -136 -352 -129 -338
rect 39 -340 47 -338
rect 83 -333 90 -317
rect 168 -332 175 -317
rect 83 -341 110 -333
rect 110 -357 118 -341
rect 168 -357 175 -340
rect -248 -370 -240 -361
rect -165 -370 -157 -361
rect 56 -370 64 -366
rect -240 -378 -236 -370
rect -228 -378 -200 -370
rect -192 -378 -157 -370
rect -148 -378 -138 -370
rect -129 -375 64 -370
rect 139 -375 147 -366
rect 186 -374 195 -277
rect 326 -340 334 -158
rect 393 -166 401 -150
rect 533 -145 540 -129
rect 533 -153 560 -145
rect 560 -169 568 -153
rect 339 -184 347 -175
rect 345 -192 351 -184
rect 359 -192 409 -184
rect 431 -188 444 -181
rect 451 -188 468 -181
rect 475 -188 490 -181
rect 506 -187 514 -178
rect 425 -203 432 -188
rect 474 -203 481 -188
rect 515 -195 518 -187
rect 526 -195 576 -187
rect 390 -229 429 -223
rect 447 -227 454 -211
rect 447 -235 474 -227
rect 474 -251 482 -235
rect 420 -268 428 -260
rect 428 -277 432 -269
rect 440 -277 460 -269
rect 468 -277 484 -269
rect 353 -294 367 -288
rect 374 -294 388 -288
rect 395 -294 440 -288
rect 448 -294 458 -288
rect 467 -294 470 -288
rect 353 -295 355 -294
rect 348 -309 355 -295
rect 397 -309 404 -294
rect 433 -309 440 -294
rect 370 -333 377 -317
rect 370 -341 397 -333
rect 397 -357 405 -341
rect 455 -357 462 -317
rect 343 -374 351 -366
rect 186 -375 351 -374
rect 426 -375 434 -366
rect 473 -375 482 -277
rect 583 -293 588 -106
rect 689 -117 696 -106
rect 738 -117 745 -102
rect 765 -108 773 -99
rect 863 -103 875 -98
rect 856 -105 875 -103
rect 882 -105 896 -98
rect 903 -105 921 -98
rect 1009 -102 1023 -95
rect 1030 -102 1044 -95
rect 1051 -102 1065 -95
rect 765 -116 777 -108
rect 785 -116 830 -108
rect 856 -120 863 -105
rect 905 -120 912 -105
rect 711 -141 718 -125
rect 1004 -117 1011 -102
rect 1053 -117 1060 -102
rect 1080 -108 1088 -99
rect 1178 -103 1190 -98
rect 1171 -105 1190 -103
rect 1197 -105 1211 -98
rect 1218 -105 1248 -98
rect 1080 -116 1092 -108
rect 1100 -116 1145 -108
rect 1171 -120 1178 -105
rect 1220 -120 1227 -105
rect 627 -153 641 -145
rect 711 -149 738 -141
rect 495 -299 504 -293
rect 510 -299 530 -293
rect 536 -299 557 -293
rect 563 -299 576 -293
rect 582 -299 588 -293
rect 495 -314 500 -299
rect 568 -314 573 -299
rect 634 -314 641 -153
rect 671 -314 679 -157
rect 738 -165 746 -149
rect 878 -144 885 -128
rect 1026 -141 1033 -125
rect 878 -152 905 -144
rect 1026 -149 1053 -141
rect 905 -168 913 -152
rect 684 -183 692 -174
rect 690 -191 696 -183
rect 704 -191 754 -183
rect 776 -187 789 -180
rect 796 -187 813 -180
rect 820 -187 835 -180
rect 851 -186 859 -177
rect 770 -202 777 -187
rect 819 -202 826 -187
rect 860 -194 863 -186
rect 871 -194 921 -186
rect 735 -228 774 -222
rect 792 -226 799 -210
rect 792 -234 819 -226
rect 819 -250 827 -234
rect 765 -267 773 -259
rect 773 -276 777 -268
rect 785 -276 805 -268
rect 813 -276 829 -268
rect 634 -322 679 -314
rect 698 -293 712 -287
rect 719 -293 733 -287
rect 740 -293 785 -287
rect 793 -293 803 -287
rect 812 -293 815 -287
rect 698 -294 700 -293
rect 693 -308 700 -294
rect 742 -308 749 -293
rect 778 -308 785 -293
rect 491 -348 497 -341
rect 541 -343 546 -323
rect 589 -338 594 -323
rect 514 -348 546 -343
rect 514 -360 520 -348
rect 589 -360 594 -344
rect 671 -339 679 -322
rect 715 -332 722 -316
rect 800 -331 807 -316
rect 715 -340 742 -332
rect 742 -356 750 -340
rect 800 -356 807 -339
rect -129 -378 68 -375
rect 56 -383 68 -378
rect 76 -383 105 -375
rect 113 -383 147 -375
rect 156 -383 166 -375
rect 175 -383 355 -375
rect 363 -383 391 -375
rect 399 -383 434 -375
rect 443 -383 453 -375
rect 462 -377 482 -375
rect 494 -377 499 -365
rect 540 -377 545 -365
rect 563 -377 569 -365
rect 688 -374 696 -365
rect 771 -374 779 -365
rect 818 -373 827 -276
rect 986 -339 994 -157
rect 1053 -165 1061 -149
rect 1193 -144 1200 -128
rect 1193 -152 1220 -144
rect 1220 -168 1228 -152
rect 999 -183 1007 -174
rect 1005 -191 1011 -183
rect 1019 -191 1069 -183
rect 1091 -187 1104 -180
rect 1111 -187 1128 -180
rect 1135 -187 1150 -180
rect 1166 -186 1174 -177
rect 1085 -202 1092 -187
rect 1134 -202 1141 -187
rect 1175 -194 1178 -186
rect 1186 -194 1236 -186
rect 1050 -228 1089 -222
rect 1107 -226 1114 -210
rect 1107 -234 1134 -226
rect 1134 -250 1142 -234
rect 1080 -267 1088 -259
rect 1088 -276 1092 -268
rect 1100 -276 1120 -268
rect 1128 -276 1144 -268
rect 1013 -293 1027 -287
rect 1034 -293 1048 -287
rect 1055 -293 1100 -287
rect 1108 -293 1118 -287
rect 1127 -293 1130 -287
rect 1013 -294 1015 -293
rect 1008 -308 1015 -294
rect 1057 -308 1064 -293
rect 1093 -308 1100 -293
rect 1030 -332 1037 -316
rect 1030 -340 1057 -332
rect 1057 -356 1065 -340
rect 1115 -356 1122 -316
rect 1003 -373 1011 -365
rect 818 -374 1011 -373
rect 1086 -374 1094 -365
rect 1133 -374 1142 -276
rect 1243 -292 1248 -105
rect 1155 -298 1164 -292
rect 1170 -298 1190 -292
rect 1196 -298 1217 -292
rect 1223 -298 1236 -292
rect 1242 -298 1248 -292
rect 1155 -313 1160 -298
rect 1228 -313 1233 -298
rect 1151 -347 1157 -340
rect 1201 -342 1206 -322
rect 1249 -338 1254 -322
rect 1174 -347 1206 -342
rect 1249 -343 1267 -338
rect 1174 -359 1180 -347
rect 1249 -359 1254 -343
rect 688 -377 700 -374
rect 462 -383 500 -377
rect 506 -383 531 -377
rect 537 -383 553 -377
rect 559 -383 572 -377
rect 578 -382 700 -377
rect 708 -382 737 -374
rect 745 -382 779 -374
rect 788 -382 798 -374
rect 807 -382 1015 -374
rect 1023 -382 1051 -374
rect 1059 -382 1094 -374
rect 1103 -382 1113 -374
rect 1122 -376 1142 -374
rect 1154 -376 1159 -364
rect 1200 -376 1205 -364
rect 1223 -376 1229 -364
rect 1122 -382 1160 -376
rect 1166 -382 1191 -376
rect 1197 -382 1213 -376
rect 1219 -382 1232 -376
rect 1238 -382 1246 -376
rect 578 -383 696 -382
rect -243 -389 -224 -383
rect -217 -389 -197 -383
rect -190 -389 -151 -383
rect -143 -389 -133 -383
rect -124 -389 -119 -383
rect -243 -404 -236 -389
rect -194 -404 -187 -389
rect -158 -404 -151 -389
rect -66 -399 98 -392
rect 385 -400 390 -397
rect -221 -428 -214 -412
rect -221 -436 -194 -428
rect -194 -452 -186 -436
rect -136 -433 -129 -412
rect 730 -415 735 -399
rect 1045 -406 1050 -393
rect 730 -422 1234 -415
rect -136 -441 -98 -433
rect -136 -452 -129 -441
rect 144 -444 157 -437
rect 164 -444 178 -437
rect 185 -444 197 -437
rect 431 -444 444 -437
rect 451 -444 465 -437
rect 472 -444 484 -437
rect 777 -444 790 -437
rect 797 -444 811 -437
rect 818 -444 830 -437
rect 1059 -444 1072 -437
rect 1079 -444 1093 -437
rect 1100 -444 1112 -437
rect 1386 -439 1399 -432
rect 1406 -439 1420 -432
rect 1427 -439 1439 -432
rect 138 -459 145 -444
rect 187 -459 194 -444
rect -248 -470 -240 -461
rect -165 -470 -157 -461
rect 425 -459 432 -444
rect 474 -459 481 -444
rect 771 -459 778 -444
rect 820 -459 827 -444
rect 1053 -459 1060 -444
rect 1102 -459 1109 -444
rect 1380 -454 1387 -439
rect 1429 -454 1436 -439
rect -240 -478 -236 -470
rect -228 -478 -200 -470
rect -192 -478 -157 -470
rect -148 -478 -138 -470
rect -129 -478 -128 -470
rect 160 -483 167 -467
rect 447 -483 454 -467
rect 793 -483 800 -467
rect 1075 -483 1082 -467
rect 1402 -478 1409 -462
rect 74 -489 137 -484
rect -243 -496 -224 -490
rect -217 -496 -198 -490
rect -190 -496 -151 -490
rect -143 -496 -133 -490
rect -124 -496 -119 -490
rect -114 -496 62 -490
rect 160 -491 187 -483
rect 207 -491 232 -483
rect 361 -489 424 -484
rect 447 -491 474 -483
rect 494 -491 519 -483
rect 707 -489 770 -484
rect 793 -491 820 -483
rect 840 -491 865 -483
rect 989 -489 1052 -484
rect 1075 -491 1102 -483
rect 1122 -491 1147 -483
rect 1316 -484 1379 -479
rect 1402 -486 1429 -478
rect 1449 -486 1474 -478
rect -243 -511 -236 -496
rect -194 -511 -187 -496
rect -158 -511 -151 -496
rect -221 -535 -214 -519
rect -136 -532 -129 -519
rect 57 -512 62 -496
rect 187 -507 195 -491
rect 474 -507 482 -491
rect 820 -507 828 -491
rect 1102 -507 1110 -491
rect 1429 -502 1437 -486
rect 62 -519 76 -512
rect 83 -519 97 -512
rect 104 -519 118 -512
rect -221 -543 -194 -535
rect -194 -559 -186 -543
rect -136 -541 -74 -532
rect 57 -534 64 -519
rect 106 -534 113 -519
rect 133 -525 141 -516
rect 231 -520 243 -515
rect 224 -522 243 -520
rect 250 -522 264 -515
rect 271 -522 289 -515
rect 349 -519 363 -512
rect 370 -519 384 -512
rect 391 -519 405 -512
rect 133 -533 145 -525
rect 153 -533 198 -525
rect -136 -559 -129 -541
rect 224 -537 231 -522
rect 273 -537 280 -522
rect 79 -558 86 -542
rect 344 -534 351 -519
rect 393 -534 400 -519
rect 420 -525 428 -516
rect 518 -520 530 -515
rect 511 -522 530 -520
rect 537 -522 551 -515
rect 558 -519 690 -515
rect 695 -519 709 -512
rect 716 -519 730 -512
rect 737 -519 751 -512
rect 558 -522 697 -519
rect 420 -533 432 -525
rect 440 -533 485 -525
rect 511 -537 518 -522
rect 560 -537 567 -522
rect 79 -566 106 -558
rect -248 -577 -240 -568
rect -165 -577 -157 -568
rect -240 -585 -236 -577
rect -228 -585 -200 -577
rect -192 -585 -157 -577
rect -148 -585 -138 -577
rect -129 -585 -128 -577
rect -243 -596 -224 -590
rect -217 -596 -198 -590
rect -190 -596 -151 -590
rect -143 -596 -133 -590
rect -124 -596 -119 -590
rect -243 -611 -236 -596
rect -194 -611 -187 -596
rect -158 -611 -151 -596
rect -259 -1052 -253 -639
rect -221 -635 -214 -619
rect -221 -643 -194 -635
rect -194 -659 -186 -643
rect -136 -637 -129 -619
rect -136 -644 -40 -637
rect -136 -659 -129 -644
rect -248 -677 -240 -668
rect -165 -677 -157 -668
rect -240 -685 -236 -677
rect -228 -685 -200 -677
rect -192 -685 -157 -677
rect -148 -685 -138 -677
rect -129 -685 -128 -677
rect -244 -711 -225 -705
rect -218 -711 -201 -705
rect -194 -711 -152 -705
rect -144 -711 -134 -705
rect -125 -711 -119 -705
rect -244 -726 -237 -711
rect -195 -726 -188 -711
rect -159 -726 -152 -711
rect -222 -750 -215 -734
rect -222 -758 -195 -750
rect -195 -774 -187 -758
rect -137 -752 -130 -734
rect 39 -738 47 -574
rect 106 -582 114 -566
rect 246 -561 253 -545
rect 366 -558 373 -542
rect 246 -569 273 -561
rect 366 -566 393 -558
rect 273 -585 281 -569
rect 52 -600 60 -591
rect 58 -608 64 -600
rect 72 -608 122 -600
rect 144 -604 157 -597
rect 164 -604 181 -597
rect 188 -604 203 -597
rect 219 -603 227 -594
rect 138 -619 145 -604
rect 187 -619 194 -604
rect 228 -611 231 -603
rect 239 -611 289 -603
rect 103 -645 142 -639
rect 160 -643 167 -627
rect 160 -651 187 -643
rect 187 -667 195 -651
rect 133 -684 141 -676
rect 141 -693 145 -685
rect 153 -693 173 -685
rect 181 -693 197 -685
rect 66 -710 80 -704
rect 87 -710 101 -704
rect 108 -710 153 -704
rect 161 -710 171 -704
rect 180 -710 183 -704
rect 66 -711 68 -710
rect 61 -725 68 -711
rect 110 -725 117 -710
rect 146 -725 153 -710
rect -78 -745 47 -738
rect -137 -759 -63 -752
rect 39 -756 47 -745
rect -137 -774 -130 -759
rect 83 -749 90 -733
rect 168 -748 175 -733
rect 83 -757 110 -749
rect 110 -773 118 -757
rect 168 -773 175 -756
rect -249 -792 -241 -783
rect -166 -792 -158 -783
rect 56 -791 64 -782
rect 139 -791 147 -782
rect 186 -790 195 -693
rect 326 -756 334 -574
rect 393 -582 401 -566
rect 533 -561 540 -545
rect 533 -569 560 -561
rect 560 -585 568 -569
rect 339 -600 347 -591
rect 345 -608 351 -600
rect 359 -608 409 -600
rect 431 -604 444 -597
rect 451 -604 468 -597
rect 475 -604 490 -597
rect 506 -603 514 -594
rect 425 -619 432 -604
rect 474 -619 481 -604
rect 515 -611 518 -603
rect 526 -611 576 -603
rect 390 -645 429 -639
rect 447 -643 454 -627
rect 447 -651 474 -643
rect 474 -667 482 -651
rect 420 -684 428 -676
rect 428 -693 432 -685
rect 440 -693 460 -685
rect 468 -693 484 -685
rect 353 -710 367 -704
rect 374 -710 388 -704
rect 395 -710 440 -704
rect 448 -710 458 -704
rect 467 -710 470 -704
rect 353 -711 355 -710
rect 348 -725 355 -711
rect 397 -725 404 -710
rect 433 -725 440 -710
rect 370 -749 377 -733
rect 370 -757 397 -749
rect 397 -773 405 -757
rect 455 -773 462 -733
rect 343 -790 351 -782
rect 186 -791 351 -790
rect 426 -791 434 -782
rect 473 -791 482 -693
rect 583 -709 588 -522
rect 690 -534 697 -522
rect 739 -534 746 -519
rect 766 -525 774 -516
rect 864 -520 876 -515
rect 857 -522 876 -520
rect 883 -522 897 -515
rect 904 -522 922 -515
rect 977 -519 991 -512
rect 998 -519 1012 -512
rect 1019 -519 1033 -512
rect 1304 -514 1318 -507
rect 1325 -514 1339 -507
rect 1346 -514 1360 -507
rect 1299 -515 1306 -514
rect 766 -533 778 -525
rect 786 -533 831 -525
rect 857 -537 864 -522
rect 906 -537 913 -522
rect 712 -558 719 -542
rect 972 -534 979 -519
rect 1021 -534 1028 -519
rect 1048 -525 1056 -516
rect 1146 -520 1158 -515
rect 1139 -522 1158 -520
rect 1165 -522 1179 -515
rect 1186 -522 1306 -515
rect 1048 -533 1060 -525
rect 1068 -533 1113 -525
rect 1139 -537 1146 -522
rect 1188 -537 1195 -522
rect 712 -566 739 -558
rect 619 -574 626 -569
rect 495 -715 504 -709
rect 510 -715 530 -709
rect 536 -715 557 -709
rect 563 -715 576 -709
rect 582 -715 588 -709
rect 495 -730 500 -715
rect 568 -730 573 -715
rect 491 -764 497 -757
rect 541 -759 546 -739
rect 589 -755 594 -739
rect 514 -764 546 -759
rect 589 -760 605 -755
rect 672 -756 680 -574
rect 739 -582 747 -566
rect 879 -561 886 -545
rect 994 -558 1001 -542
rect 879 -569 906 -561
rect 994 -566 1021 -558
rect 906 -585 914 -569
rect 685 -600 693 -591
rect 691 -608 697 -600
rect 705 -608 755 -600
rect 777 -604 790 -597
rect 797 -604 814 -597
rect 821 -604 836 -597
rect 852 -603 860 -594
rect 771 -619 778 -604
rect 820 -619 827 -604
rect 861 -611 864 -603
rect 872 -611 922 -603
rect 736 -645 775 -639
rect 793 -643 800 -627
rect 793 -651 820 -643
rect 820 -667 828 -651
rect 766 -684 774 -676
rect 774 -693 778 -685
rect 786 -693 806 -685
rect 814 -693 830 -685
rect 699 -710 713 -704
rect 720 -710 734 -704
rect 741 -710 786 -704
rect 794 -710 804 -704
rect 813 -710 816 -704
rect 699 -711 701 -710
rect 694 -725 701 -711
rect 743 -725 750 -710
rect 779 -725 786 -710
rect 514 -776 520 -764
rect 589 -776 594 -760
rect 626 -763 672 -756
rect 716 -749 723 -733
rect 801 -748 808 -733
rect 716 -757 743 -749
rect 743 -773 751 -757
rect 801 -773 808 -756
rect 56 -792 68 -791
rect -241 -800 -237 -792
rect -229 -800 -201 -792
rect -193 -800 -158 -792
rect -149 -800 -139 -792
rect -130 -799 68 -792
rect 76 -799 105 -791
rect 113 -799 147 -791
rect 156 -799 166 -791
rect 175 -799 355 -791
rect 363 -799 391 -791
rect 399 -799 434 -791
rect 443 -799 453 -791
rect 462 -793 482 -791
rect 494 -793 499 -781
rect 540 -793 545 -781
rect 563 -793 569 -781
rect 689 -791 697 -782
rect 772 -791 780 -782
rect 819 -790 828 -693
rect 954 -756 962 -574
rect 1021 -582 1029 -566
rect 1161 -561 1168 -545
rect 1161 -569 1188 -561
rect 1188 -585 1196 -569
rect 967 -600 975 -591
rect 973 -608 979 -600
rect 987 -608 1037 -600
rect 1059 -604 1072 -597
rect 1079 -604 1096 -597
rect 1103 -604 1118 -597
rect 1134 -603 1142 -594
rect 1053 -619 1060 -604
rect 1102 -619 1109 -604
rect 1143 -611 1146 -603
rect 1154 -611 1204 -603
rect 1018 -645 1057 -639
rect 1075 -643 1082 -627
rect 1075 -651 1102 -643
rect 1102 -667 1110 -651
rect 1048 -684 1056 -676
rect 1056 -693 1060 -685
rect 1068 -693 1088 -685
rect 1096 -693 1112 -685
rect 981 -710 995 -704
rect 1002 -710 1016 -704
rect 1023 -710 1068 -704
rect 1076 -710 1086 -704
rect 1095 -710 1098 -704
rect 981 -711 983 -710
rect 976 -725 983 -711
rect 1025 -725 1032 -710
rect 1061 -725 1068 -710
rect 998 -749 1005 -733
rect 998 -757 1025 -749
rect 1025 -773 1033 -757
rect 1083 -773 1090 -733
rect 971 -790 979 -782
rect 819 -791 979 -790
rect 1054 -791 1062 -782
rect 1101 -791 1110 -693
rect 1211 -709 1216 -522
rect 1299 -529 1306 -522
rect 1348 -529 1355 -514
rect 1375 -520 1383 -511
rect 1473 -515 1485 -510
rect 1466 -517 1485 -515
rect 1492 -517 1506 -510
rect 1513 -517 1531 -510
rect 1375 -528 1387 -520
rect 1395 -528 1440 -520
rect 1466 -532 1473 -517
rect 1515 -532 1522 -517
rect 1321 -553 1328 -537
rect 1321 -561 1348 -553
rect 1253 -569 1281 -561
rect 1123 -715 1132 -709
rect 1138 -715 1158 -709
rect 1164 -715 1185 -709
rect 1191 -715 1204 -709
rect 1210 -715 1216 -709
rect 1123 -730 1128 -715
rect 1196 -730 1201 -715
rect 1119 -764 1125 -757
rect 1169 -759 1174 -739
rect 1217 -754 1222 -739
rect 1281 -751 1289 -569
rect 1348 -577 1356 -561
rect 1488 -556 1495 -540
rect 1488 -564 1515 -556
rect 1515 -580 1523 -564
rect 1294 -595 1302 -586
rect 1300 -603 1306 -595
rect 1314 -603 1364 -595
rect 1386 -599 1399 -592
rect 1406 -599 1423 -592
rect 1430 -599 1445 -592
rect 1461 -598 1469 -589
rect 1380 -614 1387 -599
rect 1429 -614 1436 -599
rect 1470 -606 1473 -598
rect 1481 -606 1531 -598
rect 1345 -640 1384 -634
rect 1402 -638 1409 -622
rect 1402 -646 1429 -638
rect 1429 -662 1437 -646
rect 1375 -679 1383 -671
rect 1383 -688 1387 -680
rect 1395 -688 1415 -680
rect 1423 -688 1439 -680
rect 1308 -705 1322 -699
rect 1329 -705 1343 -699
rect 1350 -705 1395 -699
rect 1403 -705 1413 -699
rect 1422 -705 1425 -699
rect 1308 -706 1310 -705
rect 1303 -720 1310 -706
rect 1352 -720 1359 -705
rect 1388 -720 1395 -705
rect 1142 -764 1174 -759
rect 1217 -760 1234 -754
rect 1325 -744 1332 -728
rect 1410 -744 1417 -728
rect 1325 -752 1352 -744
rect 1142 -776 1148 -764
rect 1217 -776 1222 -760
rect 1352 -768 1360 -752
rect 1410 -768 1417 -751
rect 689 -793 701 -791
rect 462 -799 500 -793
rect 506 -799 531 -793
rect 537 -799 553 -793
rect 559 -799 572 -793
rect 578 -799 701 -793
rect 709 -799 738 -791
rect 746 -799 780 -791
rect 789 -799 799 -791
rect 808 -799 983 -791
rect 991 -799 1019 -791
rect 1027 -799 1062 -791
rect 1071 -799 1081 -791
rect 1090 -793 1110 -791
rect 1122 -793 1127 -781
rect 1168 -793 1173 -781
rect 1191 -793 1197 -781
rect 1298 -786 1306 -777
rect 1381 -786 1389 -777
rect 1428 -786 1437 -688
rect 1298 -793 1310 -786
rect 1090 -799 1128 -793
rect 1134 -799 1159 -793
rect 1165 -799 1181 -793
rect 1187 -799 1200 -793
rect 1206 -794 1310 -793
rect 1318 -794 1348 -786
rect 1356 -794 1389 -786
rect 1398 -794 1408 -786
rect 1417 -794 1437 -786
rect 1206 -799 1306 -794
rect -130 -800 -129 -799
rect -244 -811 -225 -805
rect -218 -811 -200 -805
rect -192 -811 -152 -805
rect -144 -811 -134 -805
rect -125 -811 -119 -805
rect 1345 -806 1581 -799
rect -244 -826 -237 -811
rect -195 -826 -188 -811
rect -159 -826 -152 -811
rect -90 -819 98 -812
rect 304 -822 385 -814
rect 731 -822 736 -816
rect 942 -820 1013 -812
rect -222 -850 -215 -834
rect -222 -858 -195 -850
rect -195 -874 -187 -858
rect -137 -851 -130 -834
rect -137 -858 -51 -851
rect -137 -874 -130 -858
rect -249 -892 -241 -883
rect -166 -892 -158 -883
rect -55 -890 731 -883
rect -241 -900 -237 -892
rect -229 -900 -201 -892
rect -193 -900 -158 -892
rect -149 -900 -139 -892
rect -130 -900 -129 -892
rect 144 -902 157 -895
rect 164 -902 178 -895
rect 185 -902 197 -895
rect 443 -902 456 -895
rect 463 -902 477 -895
rect 484 -902 496 -895
rect 758 -902 771 -895
rect 778 -902 792 -895
rect 799 -902 811 -895
rect 1087 -896 1100 -889
rect 1107 -896 1121 -889
rect 1128 -896 1140 -889
rect 1402 -896 1415 -889
rect 1422 -896 1436 -889
rect 1443 -896 1455 -889
rect -244 -918 -225 -912
rect -218 -918 -200 -912
rect -193 -918 -152 -912
rect -144 -918 -134 -912
rect -125 -918 -119 -912
rect 138 -917 145 -902
rect 187 -917 194 -902
rect -244 -933 -237 -918
rect -195 -933 -188 -918
rect -159 -933 -152 -918
rect 437 -917 444 -902
rect 486 -917 493 -902
rect 752 -917 759 -902
rect 801 -917 808 -902
rect 1081 -911 1088 -896
rect 1130 -911 1137 -896
rect 1396 -911 1403 -896
rect 1445 -911 1452 -896
rect -102 -937 94 -930
rect -222 -957 -215 -941
rect -222 -965 -195 -957
rect -195 -981 -187 -965
rect -137 -961 -130 -941
rect 160 -941 167 -925
rect 459 -941 466 -925
rect 774 -941 781 -925
rect 1103 -935 1110 -919
rect 1418 -935 1425 -919
rect 1017 -941 1080 -936
rect 71 -947 137 -942
rect 160 -949 187 -941
rect 207 -949 232 -941
rect 370 -947 436 -942
rect 459 -949 486 -941
rect 506 -949 531 -941
rect 688 -947 751 -942
rect 774 -949 801 -941
rect 821 -949 846 -941
rect 1103 -943 1130 -935
rect 1150 -943 1175 -935
rect 1332 -941 1395 -936
rect 1418 -943 1490 -935
rect -137 -968 -110 -961
rect 187 -965 195 -949
rect 486 -965 494 -949
rect 801 -965 809 -949
rect 1130 -959 1138 -943
rect 1445 -959 1453 -943
rect -137 -981 -130 -968
rect 62 -977 76 -970
rect 83 -977 100 -970
rect 107 -977 118 -970
rect -249 -999 -241 -990
rect -166 -999 -158 -990
rect 57 -992 64 -977
rect 106 -992 113 -977
rect 133 -983 141 -974
rect 231 -978 243 -973
rect 224 -980 243 -978
rect 250 -980 264 -973
rect 271 -977 356 -973
rect 361 -977 375 -970
rect 382 -977 396 -970
rect 403 -977 417 -970
rect 271 -980 363 -977
rect 133 -991 145 -983
rect 153 -991 198 -983
rect -241 -1007 -237 -999
rect -229 -1007 -201 -999
rect -193 -1007 -158 -999
rect -149 -1007 -139 -999
rect -130 -1007 -129 -999
rect 224 -995 231 -980
rect 273 -995 280 -980
rect -244 -1018 -225 -1012
rect -218 -1018 -200 -1012
rect -193 -1018 -152 -1012
rect -144 -1018 -134 -1012
rect -125 -1018 -119 -1012
rect -114 -1018 22 -1012
rect 79 -1016 86 -1000
rect 356 -992 363 -980
rect 405 -992 412 -977
rect 432 -983 440 -974
rect 530 -978 542 -973
rect 523 -980 542 -978
rect 549 -980 563 -973
rect 570 -980 588 -973
rect 676 -977 690 -970
rect 697 -977 711 -970
rect 718 -977 732 -970
rect 1005 -971 1019 -964
rect 1026 -971 1040 -964
rect 1047 -971 1061 -964
rect 910 -973 1007 -971
rect 432 -991 444 -983
rect 452 -991 497 -983
rect 523 -995 530 -980
rect 572 -995 579 -980
rect -244 -1033 -237 -1018
rect -195 -1033 -188 -1018
rect -159 -1033 -152 -1018
rect 79 -1024 106 -1016
rect -259 -1464 -253 -1058
rect -222 -1057 -215 -1041
rect -222 -1065 -195 -1057
rect -195 -1081 -187 -1065
rect -137 -1059 -130 -1041
rect -137 -1067 -93 -1059
rect -137 -1081 -130 -1067
rect -249 -1099 -241 -1090
rect -166 -1099 -158 -1090
rect -241 -1107 -237 -1099
rect -229 -1107 -201 -1099
rect -193 -1107 -158 -1099
rect -149 -1107 -139 -1099
rect -130 -1107 -129 -1099
rect -244 -1121 -225 -1115
rect -218 -1121 -202 -1115
rect -195 -1121 -152 -1115
rect -144 -1121 -134 -1115
rect -125 -1121 -119 -1115
rect -244 -1136 -237 -1121
rect -195 -1136 -188 -1121
rect -159 -1136 -152 -1121
rect -222 -1160 -215 -1144
rect -137 -1158 -130 -1144
rect -222 -1168 -195 -1160
rect -195 -1184 -187 -1168
rect -137 -1166 -7 -1158
rect -137 -1184 -130 -1166
rect 39 -1181 47 -1032
rect 106 -1040 114 -1024
rect 246 -1019 253 -1003
rect 378 -1016 385 -1000
rect 671 -992 678 -977
rect 720 -992 727 -977
rect 747 -983 755 -974
rect 845 -978 857 -973
rect 838 -980 857 -978
rect 864 -980 878 -973
rect 885 -978 1007 -973
rect 885 -980 915 -978
rect 747 -991 759 -983
rect 767 -991 812 -983
rect 838 -995 845 -980
rect 887 -995 894 -980
rect 246 -1027 273 -1019
rect 273 -1043 281 -1027
rect 52 -1058 60 -1049
rect 378 -1024 405 -1016
rect 58 -1066 64 -1058
rect 72 -1066 122 -1058
rect 144 -1062 157 -1055
rect 164 -1062 181 -1055
rect 188 -1062 203 -1055
rect 219 -1061 227 -1052
rect 138 -1077 145 -1062
rect 187 -1077 194 -1062
rect 228 -1069 231 -1061
rect 239 -1069 289 -1061
rect 103 -1103 142 -1097
rect 160 -1101 167 -1085
rect 160 -1109 187 -1101
rect 187 -1125 195 -1109
rect 133 -1142 141 -1134
rect 141 -1151 145 -1143
rect 153 -1151 173 -1143
rect 181 -1151 197 -1143
rect -67 -1187 47 -1181
rect -249 -1202 -241 -1193
rect -166 -1202 -158 -1193
rect -241 -1210 -237 -1202
rect -229 -1210 -201 -1202
rect -193 -1210 -158 -1202
rect -149 -1210 -139 -1202
rect -130 -1210 23 -1202
rect -244 -1221 -225 -1215
rect -218 -1221 -200 -1215
rect -193 -1221 -152 -1215
rect -144 -1221 -134 -1215
rect -125 -1221 -119 -1215
rect -244 -1236 -237 -1221
rect -195 -1236 -188 -1221
rect -159 -1236 -152 -1221
rect -222 -1260 -215 -1244
rect -222 -1268 -195 -1260
rect -195 -1284 -187 -1268
rect -137 -1270 -130 -1244
rect 16 -1249 23 -1210
rect 39 -1214 47 -1187
rect 66 -1168 80 -1162
rect 87 -1168 101 -1162
rect 108 -1168 153 -1162
rect 161 -1168 171 -1162
rect 180 -1168 183 -1162
rect 66 -1169 68 -1168
rect 61 -1183 68 -1169
rect 110 -1183 117 -1168
rect 146 -1183 153 -1168
rect 83 -1207 90 -1191
rect 168 -1206 175 -1191
rect 83 -1215 110 -1207
rect 110 -1231 118 -1215
rect 168 -1231 175 -1214
rect 56 -1249 64 -1240
rect 139 -1249 147 -1240
rect 186 -1248 195 -1151
rect 206 -1214 296 -1206
rect 338 -1214 346 -1027
rect 405 -1040 413 -1024
rect 545 -1019 552 -1003
rect 693 -1016 700 -1000
rect 545 -1027 572 -1019
rect 693 -1024 720 -1016
rect 572 -1043 580 -1027
rect 351 -1058 359 -1049
rect 357 -1066 363 -1058
rect 371 -1066 421 -1058
rect 443 -1062 456 -1055
rect 463 -1062 480 -1055
rect 487 -1062 502 -1055
rect 518 -1061 526 -1052
rect 437 -1077 444 -1062
rect 486 -1077 493 -1062
rect 527 -1069 530 -1061
rect 538 -1069 588 -1061
rect 402 -1103 441 -1097
rect 459 -1101 466 -1085
rect 459 -1109 486 -1101
rect 486 -1125 494 -1109
rect 432 -1142 440 -1134
rect 440 -1151 444 -1143
rect 452 -1151 472 -1143
rect 480 -1151 496 -1143
rect 365 -1168 379 -1162
rect 386 -1168 400 -1162
rect 407 -1168 452 -1162
rect 460 -1168 470 -1162
rect 479 -1168 482 -1162
rect 365 -1169 367 -1168
rect 360 -1183 367 -1169
rect 409 -1183 416 -1168
rect 445 -1183 452 -1168
rect 382 -1207 389 -1191
rect 467 -1206 474 -1191
rect 382 -1215 409 -1207
rect 409 -1231 417 -1215
rect 467 -1231 474 -1214
rect 355 -1248 363 -1240
rect 186 -1249 363 -1248
rect 438 -1249 446 -1240
rect 485 -1248 494 -1151
rect 653 -1214 661 -1032
rect 720 -1040 728 -1024
rect 860 -1019 867 -1003
rect 860 -1027 887 -1019
rect 887 -1043 895 -1027
rect 666 -1058 674 -1049
rect 672 -1066 678 -1058
rect 686 -1066 736 -1058
rect 758 -1062 771 -1055
rect 778 -1062 795 -1055
rect 802 -1062 817 -1055
rect 833 -1061 841 -1052
rect 752 -1077 759 -1062
rect 801 -1077 808 -1062
rect 842 -1069 845 -1061
rect 853 -1069 903 -1061
rect 717 -1103 756 -1097
rect 774 -1101 781 -1085
rect 774 -1109 801 -1101
rect 801 -1125 809 -1109
rect 747 -1142 755 -1134
rect 755 -1151 759 -1143
rect 767 -1151 787 -1143
rect 795 -1151 811 -1143
rect 680 -1168 694 -1162
rect 701 -1168 715 -1162
rect 722 -1168 767 -1162
rect 775 -1168 785 -1162
rect 794 -1168 797 -1162
rect 680 -1169 682 -1168
rect 675 -1183 682 -1169
rect 724 -1183 731 -1168
rect 760 -1183 767 -1168
rect 697 -1207 704 -1191
rect 697 -1215 724 -1207
rect 724 -1231 732 -1215
rect 782 -1231 789 -1191
rect 670 -1248 678 -1240
rect 485 -1249 678 -1248
rect 753 -1249 761 -1240
rect 800 -1249 809 -1151
rect 910 -1187 915 -980
rect 1000 -986 1007 -978
rect 1049 -986 1056 -971
rect 1076 -977 1084 -968
rect 1174 -972 1186 -967
rect 1167 -974 1186 -972
rect 1193 -974 1207 -967
rect 1214 -974 1232 -967
rect 1320 -971 1334 -964
rect 1341 -971 1355 -964
rect 1362 -971 1376 -964
rect 1076 -985 1088 -977
rect 1096 -985 1141 -977
rect 1167 -989 1174 -974
rect 1216 -989 1223 -974
rect 1022 -1010 1029 -994
rect 1315 -986 1322 -971
rect 1364 -986 1371 -971
rect 1391 -977 1399 -968
rect 1489 -972 1501 -967
rect 1482 -974 1501 -972
rect 1508 -974 1522 -967
rect 1529 -974 1559 -967
rect 1391 -985 1403 -977
rect 1411 -985 1456 -977
rect 1482 -989 1489 -974
rect 1531 -989 1538 -974
rect 1022 -1018 1049 -1010
rect 822 -1193 831 -1187
rect 837 -1193 857 -1187
rect 863 -1193 884 -1187
rect 890 -1193 903 -1187
rect 909 -1193 915 -1187
rect 822 -1208 827 -1193
rect 895 -1208 900 -1193
rect 954 -1208 962 -1027
rect 982 -1208 990 -1026
rect 1049 -1034 1057 -1018
rect 1189 -1013 1196 -997
rect 1337 -1010 1344 -994
rect 1189 -1021 1216 -1013
rect 1337 -1018 1364 -1010
rect 1216 -1037 1224 -1021
rect 995 -1052 1003 -1043
rect 1001 -1060 1007 -1052
rect 1015 -1060 1065 -1052
rect 1087 -1056 1100 -1049
rect 1107 -1056 1124 -1049
rect 1131 -1056 1146 -1049
rect 1162 -1055 1170 -1046
rect 1081 -1071 1088 -1056
rect 1130 -1071 1137 -1056
rect 1171 -1063 1174 -1055
rect 1182 -1063 1232 -1055
rect 1046 -1097 1085 -1091
rect 1103 -1095 1110 -1079
rect 1103 -1103 1130 -1095
rect 1130 -1119 1138 -1103
rect 1076 -1136 1084 -1128
rect 1084 -1145 1088 -1137
rect 1096 -1145 1116 -1137
rect 1124 -1145 1140 -1137
rect 1009 -1162 1023 -1156
rect 1030 -1162 1044 -1156
rect 1051 -1162 1096 -1156
rect 1104 -1162 1114 -1156
rect 1123 -1162 1126 -1156
rect 1009 -1163 1011 -1162
rect 1004 -1177 1011 -1163
rect 1053 -1177 1060 -1162
rect 1089 -1177 1096 -1162
rect 954 -1215 982 -1208
rect 1026 -1201 1033 -1185
rect 1111 -1200 1118 -1185
rect 1026 -1209 1053 -1201
rect 818 -1242 824 -1235
rect 868 -1237 873 -1217
rect 916 -1232 921 -1217
rect 1053 -1225 1061 -1209
rect 1111 -1225 1118 -1208
rect 841 -1242 873 -1237
rect 916 -1239 934 -1232
rect 16 -1257 68 -1249
rect 76 -1257 96 -1249
rect 104 -1257 147 -1249
rect 156 -1257 166 -1249
rect 175 -1257 367 -1249
rect 375 -1257 404 -1249
rect 412 -1257 446 -1249
rect 455 -1257 465 -1249
rect 474 -1257 682 -1249
rect 690 -1257 719 -1249
rect 727 -1257 761 -1249
rect 770 -1257 780 -1249
rect 789 -1257 809 -1249
rect 841 -1254 847 -1242
rect 916 -1254 921 -1239
rect -44 -1266 397 -1260
rect -137 -1277 -62 -1270
rect 144 -1276 157 -1269
rect 164 -1276 178 -1269
rect 185 -1276 197 -1269
rect 802 -1271 809 -1257
rect 821 -1271 826 -1259
rect 867 -1271 872 -1259
rect 999 -1243 1007 -1234
rect 1082 -1243 1090 -1234
rect 1129 -1242 1138 -1145
rect 1297 -1208 1305 -1026
rect 1364 -1034 1372 -1018
rect 1504 -1013 1511 -997
rect 1504 -1021 1531 -1013
rect 1531 -1037 1539 -1021
rect 1310 -1052 1318 -1043
rect 1316 -1060 1322 -1052
rect 1330 -1060 1380 -1052
rect 1402 -1056 1415 -1049
rect 1422 -1056 1439 -1049
rect 1446 -1056 1461 -1049
rect 1477 -1055 1485 -1046
rect 1396 -1071 1403 -1056
rect 1445 -1071 1452 -1056
rect 1486 -1063 1489 -1055
rect 1497 -1063 1547 -1055
rect 1361 -1097 1400 -1091
rect 1418 -1095 1425 -1079
rect 1418 -1103 1445 -1095
rect 1445 -1119 1453 -1103
rect 1391 -1136 1399 -1128
rect 1399 -1145 1403 -1137
rect 1411 -1145 1431 -1137
rect 1439 -1145 1455 -1137
rect 1324 -1162 1338 -1156
rect 1345 -1162 1359 -1156
rect 1366 -1162 1411 -1156
rect 1419 -1162 1429 -1156
rect 1438 -1162 1441 -1156
rect 1324 -1163 1326 -1162
rect 1319 -1177 1326 -1163
rect 1368 -1177 1375 -1162
rect 1404 -1177 1411 -1162
rect 1341 -1201 1348 -1185
rect 1341 -1209 1368 -1201
rect 1368 -1225 1376 -1209
rect 1426 -1225 1433 -1185
rect 1314 -1242 1322 -1234
rect 1129 -1243 1322 -1242
rect 1397 -1243 1405 -1234
rect 1444 -1243 1453 -1145
rect 1554 -1181 1559 -974
rect 1466 -1187 1475 -1181
rect 1481 -1187 1501 -1181
rect 1507 -1187 1528 -1181
rect 1534 -1187 1547 -1181
rect 1553 -1187 1559 -1181
rect 1466 -1202 1471 -1187
rect 1539 -1202 1544 -1187
rect 1462 -1236 1468 -1229
rect 1512 -1231 1517 -1211
rect 1560 -1225 1565 -1211
rect 1574 -1225 1581 -806
rect 1485 -1236 1517 -1231
rect 1560 -1232 1581 -1225
rect 999 -1251 1011 -1243
rect 1019 -1251 1048 -1243
rect 1056 -1251 1090 -1243
rect 1099 -1251 1109 -1243
rect 1118 -1251 1326 -1243
rect 1334 -1251 1362 -1243
rect 1370 -1251 1405 -1243
rect 1414 -1251 1424 -1243
rect 1433 -1251 1453 -1243
rect 1485 -1248 1491 -1236
rect 1560 -1248 1565 -1232
rect 890 -1271 896 -1259
rect 999 -1271 1007 -1251
rect -137 -1284 -130 -1277
rect 138 -1291 145 -1276
rect 187 -1291 194 -1276
rect 802 -1277 827 -1271
rect 833 -1277 858 -1271
rect 864 -1277 880 -1271
rect 886 -1277 899 -1271
rect 905 -1277 1007 -1271
rect 338 -1286 712 -1278
rect 1041 -1289 1046 -1268
rect 1446 -1265 1453 -1251
rect 1465 -1265 1470 -1253
rect 1511 -1265 1516 -1253
rect 1534 -1265 1540 -1253
rect 1446 -1271 1471 -1265
rect 1477 -1271 1502 -1265
rect 1508 -1271 1524 -1265
rect 1530 -1271 1543 -1265
rect 1549 -1271 1557 -1265
rect -249 -1302 -241 -1293
rect -166 -1302 -158 -1293
rect 303 -1298 1046 -1289
rect 1166 -1279 1356 -1274
rect -241 -1310 -237 -1302
rect -229 -1310 -201 -1302
rect -193 -1310 -158 -1302
rect -149 -1310 -139 -1302
rect -130 -1310 -129 -1302
rect -102 -1313 94 -1307
rect 160 -1315 167 -1299
rect 475 -1309 488 -1302
rect 495 -1309 509 -1302
rect 516 -1309 528 -1302
rect 790 -1309 803 -1302
rect 810 -1309 824 -1302
rect 831 -1309 843 -1302
rect 74 -1321 137 -1316
rect -244 -1328 -225 -1322
rect -218 -1328 -200 -1322
rect -193 -1328 -152 -1322
rect -144 -1328 -134 -1322
rect -125 -1328 -119 -1322
rect -114 -1328 62 -1322
rect 160 -1323 187 -1315
rect 207 -1323 232 -1315
rect -244 -1343 -237 -1328
rect -195 -1343 -188 -1328
rect -159 -1343 -152 -1328
rect -222 -1367 -215 -1351
rect -222 -1375 -195 -1367
rect -195 -1391 -187 -1375
rect -137 -1369 -130 -1351
rect 57 -1344 62 -1328
rect 187 -1339 195 -1323
rect 469 -1324 476 -1309
rect 518 -1324 525 -1309
rect 784 -1324 791 -1309
rect 833 -1324 840 -1309
rect 62 -1351 76 -1344
rect 83 -1351 101 -1344
rect 108 -1351 118 -1344
rect 57 -1366 64 -1351
rect 106 -1366 113 -1351
rect 133 -1357 141 -1348
rect 231 -1352 243 -1347
rect 224 -1354 243 -1352
rect 250 -1354 264 -1347
rect 271 -1354 393 -1347
rect 491 -1348 498 -1332
rect 806 -1348 813 -1332
rect 405 -1354 468 -1349
rect 133 -1365 145 -1357
rect 153 -1365 198 -1357
rect -137 -1376 -79 -1369
rect 224 -1369 231 -1354
rect 273 -1369 280 -1354
rect -137 -1391 -130 -1376
rect 79 -1390 86 -1374
rect 388 -1377 393 -1354
rect 491 -1356 518 -1348
rect 538 -1356 563 -1348
rect 720 -1354 783 -1349
rect 806 -1356 833 -1348
rect 853 -1356 878 -1348
rect 518 -1372 526 -1356
rect 833 -1372 841 -1356
rect 79 -1398 106 -1390
rect -249 -1409 -241 -1400
rect -166 -1409 -158 -1400
rect -33 -1406 39 -1399
rect -241 -1417 -237 -1409
rect -229 -1417 -201 -1409
rect -193 -1417 -158 -1409
rect -149 -1417 -139 -1409
rect -130 -1417 -129 -1409
rect -244 -1428 -225 -1422
rect -218 -1428 -201 -1422
rect -195 -1428 -152 -1422
rect -144 -1428 -134 -1422
rect -125 -1428 -119 -1422
rect -244 -1443 -237 -1428
rect -195 -1443 -188 -1428
rect -159 -1443 -152 -1428
rect -222 -1467 -215 -1451
rect -222 -1475 -195 -1467
rect -195 -1491 -187 -1475
rect -137 -1491 -130 -1451
rect -249 -1509 -241 -1500
rect -166 -1509 -158 -1500
rect -241 -1517 -237 -1509
rect -229 -1517 -201 -1509
rect -193 -1517 -158 -1509
rect -149 -1517 -139 -1509
rect -130 -1517 -129 -1509
rect -140 -1622 -129 -1517
rect 39 -1588 47 -1406
rect 106 -1414 114 -1398
rect 246 -1393 253 -1377
rect 393 -1384 407 -1377
rect 414 -1384 428 -1377
rect 435 -1384 449 -1377
rect 246 -1401 273 -1393
rect 281 -1401 350 -1393
rect 388 -1399 395 -1384
rect 437 -1399 444 -1384
rect 464 -1390 472 -1381
rect 562 -1385 574 -1380
rect 555 -1387 574 -1385
rect 581 -1387 595 -1380
rect 602 -1387 620 -1380
rect 708 -1384 722 -1377
rect 729 -1384 743 -1377
rect 750 -1384 764 -1377
rect 464 -1398 476 -1390
rect 484 -1398 529 -1390
rect 273 -1417 281 -1401
rect 555 -1402 562 -1387
rect 604 -1402 611 -1387
rect 52 -1432 60 -1423
rect 410 -1423 417 -1407
rect 703 -1399 710 -1384
rect 752 -1399 759 -1384
rect 779 -1390 787 -1381
rect 877 -1385 889 -1380
rect 870 -1387 889 -1385
rect 896 -1387 910 -1380
rect 917 -1387 947 -1380
rect 779 -1398 791 -1390
rect 799 -1398 844 -1390
rect 870 -1402 877 -1387
rect 919 -1402 926 -1387
rect 58 -1440 64 -1432
rect 72 -1440 122 -1432
rect 144 -1436 157 -1429
rect 164 -1436 181 -1429
rect 188 -1436 203 -1429
rect 219 -1435 227 -1426
rect 410 -1431 437 -1423
rect 138 -1451 145 -1436
rect 187 -1451 194 -1436
rect 228 -1443 231 -1435
rect 239 -1443 289 -1435
rect 103 -1477 142 -1471
rect 160 -1475 167 -1459
rect 160 -1483 187 -1475
rect 187 -1499 195 -1483
rect 133 -1516 141 -1508
rect 141 -1525 145 -1517
rect 153 -1525 173 -1517
rect 181 -1525 197 -1517
rect 66 -1542 80 -1536
rect 87 -1542 101 -1536
rect 108 -1542 153 -1536
rect 161 -1542 171 -1536
rect 180 -1542 183 -1536
rect 66 -1543 68 -1542
rect 61 -1557 68 -1543
rect 110 -1557 117 -1542
rect 146 -1557 153 -1542
rect 83 -1581 90 -1565
rect 168 -1580 175 -1565
rect 83 -1589 110 -1581
rect 110 -1605 118 -1589
rect 168 -1605 175 -1588
rect 56 -1622 64 -1614
rect -140 -1623 64 -1622
rect 139 -1623 147 -1614
rect 186 -1621 195 -1525
rect 206 -1588 330 -1580
rect 370 -1621 378 -1439
rect 437 -1447 445 -1431
rect 577 -1426 584 -1410
rect 725 -1423 732 -1407
rect 577 -1434 604 -1426
rect 725 -1431 752 -1423
rect 604 -1450 612 -1434
rect 383 -1465 391 -1456
rect 389 -1473 395 -1465
rect 403 -1473 453 -1465
rect 475 -1469 488 -1462
rect 495 -1469 512 -1462
rect 519 -1469 534 -1462
rect 550 -1468 558 -1459
rect 469 -1484 476 -1469
rect 518 -1484 525 -1469
rect 559 -1476 562 -1468
rect 570 -1476 620 -1468
rect 434 -1510 473 -1504
rect 491 -1508 498 -1492
rect 491 -1516 518 -1508
rect 518 -1532 526 -1516
rect 464 -1549 472 -1541
rect 472 -1558 476 -1550
rect 484 -1558 504 -1550
rect 512 -1558 528 -1550
rect 397 -1575 411 -1569
rect 418 -1575 432 -1569
rect 439 -1575 484 -1569
rect 492 -1575 502 -1569
rect 511 -1575 514 -1569
rect 397 -1576 399 -1575
rect 392 -1590 399 -1576
rect 441 -1590 448 -1575
rect 477 -1590 484 -1575
rect 186 -1623 345 -1621
rect -140 -1631 68 -1623
rect 76 -1631 96 -1623
rect 104 -1631 147 -1623
rect 156 -1631 166 -1623
rect 175 -1631 345 -1623
rect 356 -1628 370 -1621
rect 414 -1614 421 -1598
rect 499 -1613 506 -1598
rect 414 -1622 441 -1614
rect -140 -1996 -130 -1631
rect -55 -1642 329 -1634
rect 144 -1652 157 -1645
rect 164 -1652 178 -1645
rect 185 -1652 197 -1645
rect 138 -1667 145 -1652
rect 187 -1667 194 -1652
rect -72 -1684 94 -1679
rect 160 -1691 167 -1675
rect 321 -1677 329 -1642
rect 337 -1656 345 -1631
rect 441 -1638 449 -1622
rect 499 -1638 506 -1621
rect 387 -1656 395 -1647
rect 470 -1656 478 -1647
rect 517 -1655 526 -1558
rect 685 -1621 693 -1439
rect 752 -1447 760 -1431
rect 892 -1426 899 -1410
rect 892 -1434 919 -1426
rect 919 -1450 927 -1434
rect 698 -1465 706 -1456
rect 704 -1473 710 -1465
rect 718 -1473 768 -1465
rect 790 -1469 803 -1462
rect 810 -1469 827 -1462
rect 834 -1469 849 -1462
rect 865 -1468 873 -1459
rect 784 -1484 791 -1469
rect 833 -1484 840 -1469
rect 874 -1476 877 -1468
rect 885 -1476 935 -1468
rect 749 -1510 788 -1504
rect 806 -1508 813 -1492
rect 806 -1516 833 -1508
rect 833 -1532 841 -1516
rect 779 -1549 787 -1541
rect 787 -1558 791 -1550
rect 799 -1558 819 -1550
rect 827 -1558 843 -1550
rect 712 -1575 726 -1569
rect 733 -1575 747 -1569
rect 754 -1575 799 -1569
rect 807 -1575 817 -1569
rect 826 -1575 829 -1569
rect 712 -1576 714 -1575
rect 707 -1590 714 -1576
rect 756 -1590 763 -1575
rect 792 -1590 799 -1575
rect 729 -1614 736 -1598
rect 729 -1622 756 -1614
rect 756 -1638 764 -1622
rect 814 -1638 821 -1598
rect 702 -1655 710 -1647
rect 517 -1656 710 -1655
rect 785 -1656 793 -1647
rect 832 -1656 841 -1558
rect 942 -1594 947 -1387
rect 854 -1600 863 -1594
rect 869 -1600 889 -1594
rect 895 -1600 916 -1594
rect 922 -1600 935 -1594
rect 941 -1600 947 -1594
rect 854 -1615 859 -1600
rect 927 -1615 932 -1600
rect 850 -1649 856 -1642
rect 900 -1644 905 -1624
rect 948 -1639 953 -1624
rect 1166 -1639 1172 -1279
rect 873 -1649 905 -1644
rect 948 -1645 1172 -1639
rect 337 -1664 399 -1656
rect 407 -1664 436 -1656
rect 444 -1664 478 -1656
rect 487 -1664 497 -1656
rect 506 -1664 714 -1656
rect 722 -1664 750 -1656
rect 758 -1664 793 -1656
rect 802 -1664 812 -1656
rect 821 -1664 841 -1656
rect 873 -1661 879 -1649
rect 948 -1661 953 -1645
rect 321 -1684 429 -1677
rect 834 -1678 841 -1664
rect 853 -1678 858 -1666
rect 899 -1678 904 -1666
rect 922 -1678 928 -1666
rect 834 -1684 859 -1678
rect 865 -1684 890 -1678
rect 896 -1684 912 -1678
rect 918 -1684 931 -1678
rect 937 -1684 945 -1678
rect 74 -1697 137 -1692
rect 160 -1699 187 -1691
rect 207 -1699 232 -1691
rect 744 -1694 749 -1690
rect 187 -1715 195 -1699
rect -114 -1727 57 -1720
rect 62 -1727 76 -1720
rect 83 -1727 101 -1720
rect 108 -1727 118 -1720
rect 57 -1742 64 -1727
rect 106 -1742 113 -1727
rect 133 -1733 141 -1724
rect 231 -1728 243 -1723
rect 224 -1730 243 -1728
rect 250 -1730 264 -1723
rect 271 -1730 289 -1723
rect 133 -1741 145 -1733
rect 153 -1741 198 -1733
rect 224 -1745 231 -1730
rect 273 -1745 280 -1730
rect 79 -1766 86 -1750
rect 79 -1774 106 -1766
rect -85 -1782 39 -1775
rect 39 -1964 47 -1782
rect 106 -1790 114 -1774
rect 246 -1769 253 -1753
rect 246 -1777 273 -1769
rect 273 -1793 281 -1777
rect 52 -1808 60 -1799
rect 58 -1816 64 -1808
rect 72 -1816 122 -1808
rect 144 -1812 157 -1805
rect 164 -1812 181 -1805
rect 188 -1812 203 -1805
rect 219 -1811 227 -1802
rect 138 -1827 145 -1812
rect 187 -1827 194 -1812
rect 228 -1819 231 -1811
rect 239 -1819 289 -1811
rect 103 -1853 142 -1847
rect 160 -1851 167 -1835
rect 160 -1859 187 -1851
rect 187 -1875 195 -1859
rect 133 -1892 141 -1884
rect 141 -1901 145 -1893
rect 153 -1901 173 -1893
rect 181 -1901 197 -1893
rect 66 -1918 80 -1912
rect 87 -1918 101 -1912
rect 108 -1918 153 -1912
rect 161 -1918 171 -1912
rect 180 -1918 183 -1912
rect 66 -1919 68 -1918
rect 61 -1933 68 -1919
rect 110 -1933 117 -1918
rect 146 -1933 153 -1918
rect 83 -1957 90 -1941
rect 168 -1956 175 -1941
rect 83 -1965 110 -1957
rect 110 -1981 118 -1965
rect 168 -1981 175 -1964
rect 56 -1996 64 -1990
rect -140 -1999 64 -1996
rect 139 -1999 147 -1990
rect 186 -1999 195 -1901
rect -140 -2002 68 -1999
rect -141 -2007 68 -2002
rect 76 -2007 96 -1999
rect 104 -2007 147 -1999
rect 156 -2007 166 -1999
rect 175 -2007 195 -1999
<< m2contact >>
rect 381 386 386 391
rect 138 375 144 382
rect 197 375 203 382
rect 425 375 431 382
rect 484 375 490 382
rect 57 300 62 307
rect 118 300 124 307
rect 224 299 231 304
rect 344 300 349 307
rect 405 300 411 307
rect 198 286 203 294
rect 511 299 518 304
rect 485 286 490 294
rect -119 121 -114 127
rect 52 211 58 219
rect 138 215 144 222
rect 219 208 228 216
rect 133 126 141 135
rect 197 126 203 134
rect 61 108 66 115
rect 168 63 175 71
rect -248 32 -240 40
rect 339 211 345 219
rect 425 215 431 222
rect 506 208 515 216
rect 420 126 428 135
rect 484 126 490 134
rect 348 108 353 115
rect 485 55 491 62
rect -119 21 -114 27
rect 98 -9 103 -3
rect -74 -28 -66 -20
rect 138 -28 144 -21
rect 197 -28 203 -21
rect 425 -28 431 -21
rect 484 -28 490 -21
rect 770 -27 776 -20
rect 829 -27 835 -20
rect 1085 -27 1091 -20
rect 1144 -27 1150 -20
rect -248 -68 -240 -60
rect -119 -86 -114 -80
rect 57 -103 62 -96
rect 118 -103 124 -96
rect 224 -104 231 -99
rect 344 -103 349 -96
rect 405 -103 411 -96
rect 198 -117 203 -109
rect -86 -135 -78 -127
rect 511 -104 518 -99
rect 689 -102 694 -95
rect 750 -102 756 -95
rect 485 -117 490 -109
rect -248 -175 -240 -167
rect -119 -186 -114 -180
rect -108 -235 -102 -228
rect -248 -275 -240 -267
rect -119 -289 -114 -283
rect 52 -192 58 -184
rect 138 -188 144 -181
rect 219 -195 228 -187
rect 133 -277 141 -268
rect 197 -277 203 -269
rect 61 -295 66 -288
rect 168 -340 175 -332
rect -248 -378 -240 -370
rect 339 -192 345 -184
rect 425 -188 431 -181
rect 506 -195 515 -187
rect 420 -277 428 -268
rect 484 -277 490 -269
rect 348 -295 353 -288
rect 856 -103 863 -98
rect 1004 -102 1009 -95
rect 1065 -102 1071 -95
rect 830 -116 835 -108
rect 1171 -103 1178 -98
rect 1145 -116 1150 -108
rect 684 -191 690 -183
rect 770 -187 776 -180
rect 851 -194 860 -186
rect 765 -276 773 -267
rect 829 -276 835 -268
rect 693 -294 698 -287
rect 485 -348 491 -341
rect 589 -344 594 -338
rect 800 -339 807 -331
rect 999 -191 1005 -183
rect 1085 -187 1091 -180
rect 1166 -194 1175 -186
rect 1080 -276 1088 -267
rect 1144 -276 1150 -268
rect 1008 -294 1013 -287
rect 1145 -347 1151 -340
rect 1267 -343 1273 -338
rect -119 -389 -114 -383
rect -74 -399 -66 -392
rect 385 -405 390 -400
rect 1045 -412 1050 -406
rect 1234 -422 1241 -415
rect -98 -441 -90 -433
rect 138 -444 144 -437
rect 197 -444 203 -437
rect 425 -444 431 -437
rect 484 -444 490 -437
rect 771 -444 777 -437
rect 830 -444 836 -437
rect 1053 -444 1059 -437
rect 1112 -444 1118 -437
rect 1380 -439 1386 -432
rect 1439 -439 1445 -432
rect -248 -478 -240 -470
rect -119 -496 -114 -490
rect 57 -519 62 -512
rect 118 -519 124 -512
rect -74 -541 -67 -532
rect 224 -520 231 -515
rect 344 -519 349 -512
rect 405 -519 411 -512
rect 198 -533 203 -525
rect 511 -520 518 -515
rect 690 -519 695 -512
rect 751 -519 757 -512
rect 485 -533 490 -525
rect -248 -585 -240 -577
rect -119 -596 -114 -590
rect -40 -644 -33 -637
rect -248 -685 -240 -677
rect -119 -711 -114 -705
rect 52 -608 58 -600
rect 138 -604 144 -597
rect 219 -611 228 -603
rect 133 -693 141 -684
rect 197 -693 203 -685
rect 61 -711 66 -704
rect -86 -745 -78 -738
rect -63 -759 -55 -752
rect 168 -756 175 -748
rect 339 -608 345 -600
rect 425 -604 431 -597
rect 506 -611 515 -603
rect 420 -693 428 -684
rect 484 -693 490 -685
rect 348 -711 353 -704
rect 857 -520 864 -515
rect 972 -519 977 -512
rect 1033 -519 1039 -512
rect 1299 -514 1304 -507
rect 1360 -514 1366 -507
rect 831 -533 836 -525
rect 1139 -520 1146 -515
rect 1113 -533 1118 -525
rect 619 -580 626 -574
rect 485 -764 491 -757
rect 605 -760 611 -755
rect 685 -608 691 -600
rect 771 -604 777 -597
rect 852 -611 861 -603
rect 766 -693 774 -684
rect 830 -693 836 -685
rect 694 -711 699 -704
rect 619 -763 626 -756
rect 801 -756 808 -748
rect -249 -800 -241 -792
rect 967 -608 973 -600
rect 1053 -604 1059 -597
rect 1134 -611 1143 -603
rect 1048 -693 1056 -684
rect 1112 -693 1118 -685
rect 976 -711 981 -704
rect 1466 -515 1473 -510
rect 1440 -528 1445 -520
rect 1113 -764 1119 -757
rect 1294 -603 1300 -595
rect 1380 -599 1386 -592
rect 1461 -606 1470 -598
rect 1375 -688 1383 -679
rect 1439 -688 1445 -680
rect 1303 -706 1308 -699
rect 1234 -760 1241 -754
rect 1410 -751 1417 -744
rect -119 -811 -114 -805
rect -98 -819 -90 -812
rect 296 -822 304 -814
rect 934 -820 942 -812
rect 731 -828 736 -822
rect -51 -858 -44 -851
rect -63 -890 -55 -883
rect 731 -890 736 -883
rect -249 -900 -241 -892
rect 138 -902 144 -895
rect 197 -902 203 -895
rect 437 -902 443 -895
rect 496 -902 502 -895
rect 752 -902 758 -895
rect 811 -902 817 -895
rect 1081 -896 1087 -889
rect 1140 -896 1146 -889
rect 1396 -896 1402 -889
rect 1455 -896 1461 -889
rect -119 -918 -114 -912
rect -108 -937 -102 -930
rect -110 -968 -102 -961
rect 57 -977 62 -970
rect 118 -977 124 -970
rect 224 -978 231 -973
rect 356 -977 361 -970
rect 417 -977 423 -970
rect 198 -991 203 -983
rect -249 -1007 -241 -999
rect -119 -1018 -114 -1012
rect 22 -1018 27 -1012
rect 523 -978 530 -973
rect 671 -977 676 -970
rect 732 -977 738 -970
rect 1000 -971 1005 -964
rect 1061 -971 1067 -964
rect 497 -991 502 -983
rect -93 -1067 -85 -1059
rect -249 -1107 -241 -1099
rect -119 -1121 -114 -1115
rect -7 -1166 1 -1158
rect 838 -978 845 -973
rect 812 -991 817 -983
rect 52 -1066 58 -1058
rect 138 -1062 144 -1055
rect 219 -1069 228 -1061
rect 133 -1151 141 -1142
rect 197 -1151 203 -1143
rect -74 -1187 -67 -1181
rect -249 -1210 -241 -1202
rect -119 -1221 -114 -1215
rect 61 -1169 66 -1162
rect 168 -1214 175 -1206
rect 199 -1214 206 -1206
rect 296 -1214 304 -1206
rect 351 -1066 357 -1058
rect 437 -1062 443 -1055
rect 518 -1069 527 -1061
rect 432 -1151 440 -1142
rect 496 -1151 502 -1143
rect 360 -1169 365 -1162
rect 467 -1214 474 -1206
rect 666 -1066 672 -1058
rect 752 -1062 758 -1055
rect 833 -1069 842 -1061
rect 747 -1151 755 -1142
rect 811 -1151 817 -1143
rect 675 -1169 680 -1162
rect 1167 -972 1174 -967
rect 1315 -971 1320 -964
rect 1376 -971 1382 -964
rect 1141 -985 1146 -977
rect 1482 -972 1489 -967
rect 1456 -985 1461 -977
rect 995 -1060 1001 -1052
rect 1081 -1056 1087 -1049
rect 1162 -1063 1171 -1055
rect 1076 -1145 1084 -1136
rect 1140 -1145 1146 -1137
rect 1004 -1163 1009 -1156
rect 812 -1242 818 -1235
rect 1111 -1208 1118 -1200
rect 934 -1239 942 -1232
rect -51 -1266 -44 -1260
rect -62 -1277 -55 -1270
rect 138 -1276 144 -1269
rect 197 -1276 203 -1269
rect 1310 -1060 1316 -1052
rect 1396 -1056 1402 -1049
rect 1477 -1063 1486 -1055
rect 1391 -1145 1399 -1136
rect 1455 -1145 1461 -1137
rect 1319 -1163 1324 -1156
rect 1456 -1236 1462 -1229
rect 330 -1286 338 -1278
rect 295 -1298 303 -1289
rect -249 -1310 -241 -1302
rect -110 -1313 -102 -1307
rect 469 -1309 475 -1302
rect 528 -1309 534 -1302
rect 784 -1309 790 -1302
rect 843 -1309 849 -1302
rect -119 -1328 -114 -1322
rect 57 -1351 62 -1344
rect 118 -1351 124 -1344
rect 224 -1352 231 -1347
rect 198 -1365 203 -1357
rect -79 -1376 -72 -1369
rect -40 -1406 -33 -1399
rect -249 -1417 -241 -1409
rect -119 -1428 -114 -1422
rect -249 -1517 -241 -1509
rect 388 -1384 393 -1377
rect 449 -1384 455 -1377
rect 350 -1401 356 -1393
rect 555 -1385 562 -1380
rect 703 -1384 708 -1377
rect 764 -1384 770 -1377
rect 529 -1398 534 -1390
rect 870 -1385 877 -1380
rect 844 -1398 849 -1390
rect 52 -1440 58 -1432
rect 138 -1436 144 -1429
rect 219 -1443 228 -1435
rect 133 -1525 141 -1516
rect 197 -1525 203 -1517
rect 61 -1543 66 -1536
rect 168 -1588 175 -1580
rect 199 -1588 206 -1580
rect 330 -1588 338 -1580
rect 383 -1473 389 -1465
rect 469 -1469 475 -1462
rect 550 -1476 559 -1468
rect 464 -1558 472 -1549
rect 528 -1558 534 -1550
rect 392 -1576 397 -1569
rect 350 -1628 356 -1621
rect -62 -1642 -55 -1634
rect 138 -1652 144 -1645
rect 197 -1652 203 -1645
rect -79 -1684 -72 -1679
rect 499 -1621 506 -1613
rect 698 -1473 704 -1465
rect 784 -1469 790 -1462
rect 865 -1476 874 -1468
rect 779 -1558 787 -1549
rect 843 -1558 849 -1550
rect 707 -1576 712 -1569
rect 844 -1649 850 -1642
rect 744 -1699 749 -1694
rect -119 -1727 -114 -1720
rect 57 -1727 62 -1720
rect 118 -1727 124 -1720
rect 224 -1728 231 -1723
rect 198 -1741 203 -1733
rect -93 -1782 -85 -1775
rect 52 -1816 58 -1808
rect 138 -1812 144 -1805
rect 219 -1819 228 -1811
rect 133 -1901 141 -1892
rect 197 -1901 203 -1893
rect 61 -1919 66 -1912
rect 168 -1964 175 -1956
<< metal2 >>
rect 386 386 620 391
rect 125 375 138 382
rect 203 375 425 382
rect 490 375 518 382
rect 125 307 132 375
rect 29 300 57 307
rect 124 300 132 307
rect 29 127 35 300
rect 125 222 132 300
rect 224 374 419 375
rect 224 304 231 374
rect 412 307 419 374
rect 317 300 344 307
rect 411 300 419 307
rect 198 234 203 286
rect 198 227 215 234
rect -114 121 35 127
rect 125 215 138 222
rect 209 216 215 227
rect 52 135 58 211
rect 209 208 219 216
rect 52 126 133 135
rect 219 134 228 208
rect 203 126 228 134
rect -294 32 -248 40
rect -294 -60 -286 32
rect -118 27 -114 121
rect 29 115 35 121
rect 317 115 322 300
rect 412 222 419 300
rect 511 304 518 375
rect 485 234 490 286
rect 485 227 502 234
rect 412 215 425 222
rect 496 216 502 227
rect 339 135 345 211
rect 496 208 506 216
rect 339 126 420 135
rect 506 134 515 208
rect 490 126 515 134
rect 29 108 61 115
rect 317 108 348 115
rect 175 63 287 71
rect -294 -68 -248 -60
rect -294 -167 -286 -68
rect -118 -80 -114 21
rect 279 16 287 63
rect 471 55 485 62
rect 471 16 477 55
rect 279 9 477 16
rect 103 -9 609 -3
rect -294 -175 -248 -167
rect -294 -267 -286 -175
rect -118 -180 -114 -86
rect -294 -275 -248 -267
rect -294 -370 -286 -275
rect -118 -283 -114 -186
rect -294 -378 -248 -370
rect -294 -470 -286 -378
rect -118 -383 -114 -289
rect -294 -478 -248 -470
rect -294 -577 -286 -478
rect -118 -490 -114 -389
rect -108 -433 -102 -235
rect -110 -441 -102 -433
rect -294 -585 -248 -577
rect -294 -677 -286 -585
rect -118 -590 -114 -496
rect -294 -685 -248 -677
rect -294 -792 -286 -685
rect -118 -705 -114 -596
rect -294 -800 -249 -792
rect -294 -892 -286 -800
rect -118 -805 -114 -711
rect -294 -900 -249 -892
rect -294 -999 -286 -900
rect -118 -912 -114 -811
rect -294 -1007 -249 -999
rect -294 -1099 -286 -1007
rect -118 -1012 -114 -918
rect -108 -930 -102 -441
rect -98 -812 -90 -441
rect -86 -738 -78 -135
rect -74 -392 -66 -28
rect 125 -28 138 -21
rect 203 -28 425 -21
rect 490 -28 518 -21
rect 125 -96 132 -28
rect 29 -103 57 -96
rect 124 -103 132 -96
rect 29 -288 35 -103
rect 125 -181 132 -103
rect 224 -29 419 -28
rect 224 -99 231 -29
rect 412 -96 419 -29
rect 317 -103 344 -96
rect 411 -103 419 -96
rect 198 -169 203 -117
rect 198 -176 215 -169
rect 125 -188 138 -181
rect 209 -187 215 -176
rect 52 -268 58 -192
rect 209 -195 219 -187
rect 52 -277 133 -268
rect 219 -269 228 -195
rect 203 -277 228 -269
rect 317 -288 322 -103
rect 412 -181 419 -103
rect 511 -99 518 -28
rect 485 -169 490 -117
rect 485 -176 502 -169
rect 412 -188 425 -181
rect 496 -187 502 -176
rect 339 -268 345 -192
rect 496 -195 506 -187
rect 339 -277 420 -268
rect 506 -269 515 -195
rect 490 -277 515 -269
rect 29 -295 61 -288
rect 317 -295 348 -288
rect 175 -340 287 -332
rect 602 -338 609 -9
rect 613 -7 620 386
rect 613 -14 1273 -7
rect 757 -27 770 -20
rect 835 -27 1085 -20
rect 1150 -27 1178 -20
rect 757 -95 764 -27
rect 661 -102 689 -95
rect 756 -102 764 -95
rect 661 -287 667 -102
rect 757 -180 764 -102
rect 856 -28 1079 -27
rect 856 -98 863 -28
rect 1072 -95 1079 -28
rect 977 -102 1004 -95
rect 1071 -102 1079 -95
rect 830 -168 835 -116
rect 830 -175 847 -168
rect 757 -187 770 -180
rect 841 -186 847 -175
rect 684 -267 690 -191
rect 841 -194 851 -186
rect 684 -276 765 -267
rect 851 -268 860 -194
rect 835 -276 860 -268
rect 977 -287 982 -102
rect 1072 -180 1079 -102
rect 1171 -98 1178 -27
rect 1145 -168 1150 -116
rect 1145 -175 1162 -168
rect 1072 -187 1085 -180
rect 1156 -186 1162 -175
rect 999 -267 1005 -191
rect 1156 -194 1166 -186
rect 999 -276 1080 -267
rect 1166 -268 1175 -194
rect 1150 -276 1175 -268
rect 661 -294 693 -287
rect 977 -294 1008 -287
rect 279 -387 287 -340
rect 469 -348 485 -341
rect 594 -344 609 -338
rect 807 -339 919 -331
rect 469 -387 473 -348
rect 279 -392 473 -387
rect 477 -374 612 -370
rect 477 -401 480 -374
rect 390 -405 480 -401
rect 125 -444 138 -437
rect 203 -444 425 -437
rect 490 -444 518 -437
rect 125 -512 132 -444
rect 29 -519 57 -512
rect 124 -519 132 -512
rect -294 -1107 -249 -1099
rect -294 -1202 -286 -1107
rect -118 -1115 -114 -1018
rect -294 -1210 -249 -1202
rect -294 -1302 -286 -1210
rect -118 -1215 -114 -1121
rect -294 -1310 -249 -1302
rect -294 -1409 -286 -1310
rect -118 -1322 -114 -1221
rect -110 -1307 -102 -968
rect -294 -1417 -249 -1409
rect -294 -1509 -286 -1417
rect -118 -1422 -114 -1328
rect -294 -1517 -249 -1509
rect -119 -1720 -114 -1428
rect -93 -1775 -85 -1067
rect -74 -1181 -67 -541
rect -63 -883 -55 -759
rect -51 -1260 -44 -858
rect -79 -1679 -72 -1376
rect -62 -1634 -55 -1277
rect -40 -1399 -33 -644
rect 29 -704 35 -519
rect 125 -597 132 -519
rect 224 -445 419 -444
rect 224 -515 231 -445
rect 412 -512 419 -445
rect 317 -519 344 -512
rect 411 -519 419 -512
rect 198 -585 203 -533
rect 198 -592 215 -585
rect 125 -604 138 -597
rect 209 -603 215 -592
rect 52 -684 58 -608
rect 209 -611 219 -603
rect 52 -693 133 -684
rect 219 -685 228 -611
rect 203 -693 228 -685
rect 317 -704 322 -519
rect 412 -597 419 -519
rect 511 -515 518 -444
rect 605 -438 612 -374
rect 911 -395 919 -339
rect 1267 -338 1273 -14
rect 1127 -347 1145 -340
rect 1127 -395 1132 -347
rect 911 -402 1132 -395
rect 1136 -375 1546 -369
rect 1136 -406 1141 -375
rect 1050 -412 1141 -406
rect 485 -585 490 -533
rect 485 -592 502 -585
rect 412 -604 425 -597
rect 496 -603 502 -592
rect 339 -684 345 -608
rect 496 -611 506 -603
rect 339 -693 420 -684
rect 506 -685 515 -611
rect 490 -693 515 -685
rect 29 -711 61 -704
rect 317 -711 348 -704
rect 175 -756 287 -748
rect 279 -803 287 -756
rect 605 -755 611 -438
rect 758 -444 771 -437
rect 836 -444 1053 -437
rect 1118 -444 1146 -437
rect 758 -512 765 -444
rect 662 -519 690 -512
rect 757 -519 765 -512
rect 475 -764 485 -757
rect 619 -756 626 -580
rect 662 -704 668 -519
rect 758 -597 765 -519
rect 857 -445 1047 -444
rect 857 -515 864 -445
rect 1040 -512 1047 -445
rect 945 -519 972 -512
rect 1039 -519 1047 -512
rect 831 -585 836 -533
rect 831 -592 848 -585
rect 758 -604 771 -597
rect 842 -603 848 -592
rect 685 -684 691 -608
rect 842 -611 852 -603
rect 685 -693 766 -684
rect 852 -685 861 -611
rect 836 -693 861 -685
rect 945 -704 950 -519
rect 1040 -597 1047 -519
rect 1139 -515 1146 -444
rect 1113 -585 1118 -533
rect 1113 -592 1130 -585
rect 1040 -604 1053 -597
rect 1124 -603 1130 -592
rect 967 -684 973 -608
rect 1124 -611 1134 -603
rect 967 -693 1048 -684
rect 1134 -685 1143 -611
rect 1118 -693 1143 -685
rect 662 -711 694 -704
rect 945 -711 976 -704
rect 808 -756 920 -748
rect 475 -803 482 -764
rect 279 -810 482 -803
rect 912 -801 920 -756
rect 1234 -754 1241 -422
rect 1367 -439 1380 -432
rect 1445 -439 1473 -432
rect 1367 -507 1374 -439
rect 1269 -514 1299 -507
rect 1366 -514 1374 -507
rect 1269 -699 1277 -514
rect 1367 -592 1374 -514
rect 1466 -510 1473 -439
rect 1440 -580 1445 -528
rect 1440 -587 1457 -580
rect 1367 -599 1380 -592
rect 1451 -598 1457 -587
rect 1294 -679 1300 -603
rect 1451 -606 1461 -598
rect 1294 -688 1375 -679
rect 1461 -680 1470 -606
rect 1445 -688 1470 -680
rect 1269 -706 1303 -699
rect 1538 -744 1546 -375
rect 1417 -751 1546 -744
rect 1102 -764 1113 -757
rect 1102 -801 1109 -764
rect 912 -808 1109 -801
rect 125 -902 138 -895
rect 203 -902 231 -895
rect 125 -970 132 -902
rect 27 -977 57 -970
rect 124 -977 132 -970
rect -7 -1634 1 -1166
rect 27 -1162 35 -977
rect 125 -1055 132 -977
rect 224 -973 231 -902
rect 198 -1043 203 -991
rect 198 -1050 215 -1043
rect 125 -1062 138 -1055
rect 209 -1061 215 -1050
rect 52 -1142 58 -1066
rect 209 -1069 219 -1061
rect 52 -1151 133 -1142
rect 219 -1143 228 -1069
rect 203 -1151 228 -1143
rect 27 -1169 61 -1162
rect 296 -1206 304 -822
rect 731 -883 736 -828
rect 424 -902 437 -895
rect 502 -902 752 -895
rect 817 -902 845 -895
rect 424 -970 431 -902
rect 328 -977 356 -970
rect 423 -977 431 -970
rect 328 -1162 334 -977
rect 424 -1055 431 -977
rect 523 -903 746 -902
rect 523 -973 530 -903
rect 739 -970 746 -903
rect 644 -977 671 -970
rect 738 -977 746 -970
rect 497 -1043 502 -991
rect 497 -1050 514 -1043
rect 424 -1062 437 -1055
rect 508 -1061 514 -1050
rect 351 -1142 357 -1066
rect 508 -1069 518 -1061
rect 351 -1151 432 -1142
rect 518 -1143 527 -1069
rect 502 -1151 527 -1143
rect 644 -1162 649 -977
rect 739 -1055 746 -977
rect 838 -973 845 -902
rect 812 -1043 817 -991
rect 812 -1050 829 -1043
rect 739 -1062 752 -1055
rect 823 -1061 829 -1050
rect 666 -1142 672 -1066
rect 823 -1069 833 -1061
rect 666 -1151 747 -1142
rect 833 -1143 842 -1069
rect 817 -1151 842 -1143
rect 328 -1169 360 -1162
rect 644 -1169 675 -1162
rect 175 -1214 199 -1206
rect 474 -1214 586 -1206
rect 125 -1276 138 -1269
rect 203 -1276 231 -1269
rect 125 -1344 132 -1276
rect 27 -1351 57 -1344
rect 124 -1351 132 -1344
rect 27 -1536 35 -1351
rect 125 -1429 132 -1351
rect 224 -1347 231 -1276
rect 578 -1270 586 -1214
rect 934 -1232 942 -820
rect 1068 -896 1081 -889
rect 1146 -896 1396 -889
rect 1461 -896 1489 -889
rect 1068 -964 1075 -896
rect 972 -971 1000 -964
rect 1067 -971 1075 -964
rect 972 -1156 978 -971
rect 1068 -1049 1075 -971
rect 1167 -897 1390 -896
rect 1167 -967 1174 -897
rect 1383 -964 1390 -897
rect 1288 -971 1315 -964
rect 1382 -971 1390 -964
rect 1141 -1037 1146 -985
rect 1141 -1044 1158 -1037
rect 1068 -1056 1081 -1049
rect 1152 -1055 1158 -1044
rect 995 -1136 1001 -1060
rect 1152 -1063 1162 -1055
rect 995 -1145 1076 -1136
rect 1162 -1137 1171 -1063
rect 1146 -1145 1171 -1137
rect 1288 -1156 1293 -971
rect 1383 -1049 1390 -971
rect 1482 -967 1489 -896
rect 1456 -1037 1461 -985
rect 1456 -1044 1473 -1037
rect 1383 -1056 1396 -1049
rect 1467 -1055 1473 -1044
rect 1310 -1136 1316 -1060
rect 1467 -1063 1477 -1055
rect 1310 -1145 1391 -1136
rect 1477 -1137 1486 -1063
rect 1461 -1145 1486 -1137
rect 972 -1163 1004 -1156
rect 1288 -1163 1319 -1156
rect 1118 -1208 1230 -1200
rect 804 -1242 812 -1235
rect 804 -1270 809 -1242
rect 578 -1277 809 -1270
rect 1222 -1264 1230 -1208
rect 1448 -1236 1456 -1229
rect 1448 -1264 1453 -1236
rect 1222 -1271 1453 -1264
rect 198 -1417 203 -1365
rect 198 -1424 215 -1417
rect 125 -1436 138 -1429
rect 209 -1435 215 -1424
rect 52 -1516 58 -1440
rect 209 -1443 219 -1435
rect 52 -1525 133 -1516
rect 219 -1517 228 -1443
rect 203 -1525 228 -1517
rect 27 -1543 61 -1536
rect 175 -1588 199 -1580
rect 295 -1634 303 -1298
rect 330 -1580 338 -1286
rect 456 -1309 469 -1302
rect 534 -1309 784 -1302
rect 849 -1309 877 -1302
rect 456 -1377 463 -1309
rect 360 -1384 388 -1377
rect 455 -1384 463 -1377
rect 350 -1621 356 -1401
rect 360 -1569 366 -1384
rect 456 -1462 463 -1384
rect 555 -1310 778 -1309
rect 555 -1380 562 -1310
rect 771 -1377 778 -1310
rect 676 -1384 703 -1377
rect 770 -1384 778 -1377
rect 529 -1450 534 -1398
rect 529 -1457 546 -1450
rect 456 -1469 469 -1462
rect 540 -1468 546 -1457
rect 383 -1549 389 -1473
rect 540 -1476 550 -1468
rect 383 -1558 464 -1549
rect 550 -1550 559 -1476
rect 534 -1558 559 -1550
rect 676 -1569 681 -1384
rect 771 -1462 778 -1384
rect 870 -1380 877 -1309
rect 844 -1450 849 -1398
rect 844 -1457 861 -1450
rect 771 -1469 784 -1462
rect 855 -1468 861 -1457
rect 698 -1549 704 -1473
rect 855 -1476 865 -1468
rect 698 -1558 779 -1549
rect 865 -1550 874 -1476
rect 849 -1558 874 -1550
rect 360 -1576 392 -1569
rect 676 -1576 707 -1569
rect 506 -1621 618 -1613
rect -7 -1640 303 -1634
rect 125 -1652 138 -1645
rect 203 -1652 231 -1645
rect 125 -1720 132 -1652
rect 27 -1727 57 -1720
rect 124 -1727 132 -1720
rect 27 -1912 35 -1727
rect 125 -1805 132 -1727
rect 224 -1723 231 -1652
rect 610 -1677 618 -1621
rect 836 -1649 844 -1642
rect 836 -1677 841 -1649
rect 610 -1684 841 -1677
rect 198 -1793 203 -1741
rect 198 -1800 215 -1793
rect 125 -1812 138 -1805
rect 209 -1811 215 -1800
rect 52 -1892 58 -1816
rect 209 -1819 219 -1811
rect 52 -1901 133 -1892
rect 219 -1893 228 -1819
rect 203 -1901 228 -1893
rect 27 -1919 61 -1912
rect 744 -1956 749 -1699
rect 175 -1964 749 -1956
<< labels >>
rlabel metal1 -243 121 -122 127 5 drain
rlabel metal1 -248 -68 -157 -60 1 Gnd
rlabel metal1 -243 21 -122 27 5 drain
rlabel metal1 -248 -175 -157 -167 1 Gnd
rlabel metal1 -243 -86 -122 -80 5 drain
rlabel metal1 -243 -186 -122 -180 5 drain
rlabel metal1 -243 -596 -122 -590 5 drain
rlabel metal1 -248 -685 -157 -677 1 Gnd
rlabel metal1 -243 -496 -122 -490 5 drain
rlabel metal1 -248 -585 -157 -577 1 Gnd
rlabel metal1 -243 -389 -122 -383 5 drain
rlabel metal1 -248 -478 -157 -470 1 Gnd
rlabel metal1 -248 -378 -157 -370 1 Gnd
rlabel metal1 -249 -1210 -158 -1202 1 Gnd
rlabel metal1 -244 -1121 -123 -1115 5 drain
rlabel metal1 -249 -1310 -158 -1302 1 Gnd
rlabel metal1 -244 -1221 -123 -1215 5 drain
rlabel metal1 -249 -1417 -158 -1409 1 Gnd
rlabel metal1 -244 -1328 -123 -1322 5 drain
rlabel metal1 -249 -1517 -158 -1509 1 Gnd
rlabel metal1 -244 -1428 -123 -1422 5 drain
rlabel metal1 -244 -1018 -123 -1012 5 drain
rlabel metal1 -249 -1107 -158 -1099 1 Gnd
rlabel metal1 -244 -918 -123 -912 5 drain
rlabel metal1 -249 -1007 -158 -999 1 Gnd
rlabel metal1 -244 -811 -123 -805 5 drain
rlabel metal1 -249 -900 -158 -892 1 Gnd
rlabel metal1 -244 -711 -123 -705 5 drain
rlabel metal1 -249 -800 -158 -792 1 Gnd
rlabel metal1 -248 32 -157 40 1 Gnd
rlabel metal1 -243 -289 -122 -283 5 drain
rlabel metal1 -248 -275 -157 -267 1 Gnd
rlabel polysilicon -206 -38 -201 -30 1 A3
rlabel polysilicon -206 -449 -201 -441 1 A2
rlabel polysilicon -207 -871 -202 -863 1 A1
rlabel polysilicon -207 -1281 -202 -1273 1 A0
rlabel polysilicon -234 67 -229 75 1 B3
rlabel polysilicon -234 -35 -229 -27 1 B2
rlabel polysilicon -234 -139 -229 -131 1 B1
rlabel polysilicon -234 -236 -229 -228 1 B0
rlabel metal1 -137 -1478 -130 -1466 1 P0
rlabel metal1 57 -977 122 -970 5 drain
rlabel metal1 52 -1066 122 -1058 1 Gnd
rlabel metal1 219 -1069 289 -1061 1 Gnd
rlabel metal1 224 -980 289 -973 5 drain
rlabel metal1 57 -1351 122 -1344 5 drain
rlabel metal1 52 -1440 122 -1432 1 Gnd
rlabel metal1 219 -1443 289 -1435 1 Gnd
rlabel metal1 224 -1354 289 -1347 5 drain
rlabel metal1 224 297 289 304 5 drain
rlabel metal1 219 208 289 216 1 Gnd
rlabel metal1 52 211 122 219 1 Gnd
rlabel metal1 57 300 122 307 5 drain
rlabel metal1 511 297 576 304 5 drain
rlabel metal1 506 208 576 216 1 Gnd
rlabel metal1 339 211 409 219 1 Gnd
rlabel metal1 344 300 409 307 5 drain
rlabel metal1 560 234 568 258 1 P6
rlabel metal1 589 58 594 66 1 C5
rlabel metal1 57 -103 122 -96 5 drain
rlabel metal1 52 -192 122 -184 1 Gnd
rlabel metal1 219 -195 289 -187 1 Gnd
rlabel metal1 224 -106 289 -99 5 drain
rlabel metal1 344 -103 409 -96 5 drain
rlabel metal1 339 -192 409 -184 1 Gnd
rlabel metal1 506 -195 576 -187 1 Gnd
rlabel metal1 511 -106 576 -99 5 drain
rlabel metal1 856 -105 921 -98 5 drain
rlabel metal1 851 -194 921 -186 1 Gnd
rlabel metal1 684 -191 754 -183 1 Gnd
rlabel metal1 689 -102 754 -95 5 drain
rlabel metal1 1171 -105 1236 -98 5 drain
rlabel metal1 1166 -194 1236 -186 1 Gnd
rlabel metal1 999 -191 1069 -183 1 Gnd
rlabel metal1 1004 -102 1069 -95 5 drain
rlabel metal1 1220 -168 1228 -144 1 P5
rlabel metal1 857 -522 922 -515 5 drain
rlabel metal1 852 -611 922 -603 1 Gnd
rlabel metal1 685 -608 755 -600 1 Gnd
rlabel metal1 972 -519 1037 -512 5 drain
rlabel metal1 967 -608 1037 -600 1 Gnd
rlabel metal1 1134 -611 1204 -603 1 Gnd
rlabel metal1 1139 -522 1204 -515 5 drain
rlabel metal1 1515 -580 1523 -556 1 P4
rlabel metal1 1299 -514 1364 -507 5 drain
rlabel metal1 1294 -603 1364 -595 1 Gnd
rlabel metal1 1461 -606 1531 -598 1 Gnd
rlabel metal1 1466 -517 1531 -510 5 drain
rlabel metal1 57 -519 122 -512 5 drain
rlabel metal1 52 -608 122 -600 1 Gnd
rlabel metal1 219 -611 289 -603 1 Gnd
rlabel metal1 224 -522 289 -515 5 drain
rlabel metal1 344 -519 409 -512 5 drain
rlabel metal1 339 -608 409 -600 1 Gnd
rlabel metal1 506 -611 576 -603 1 Gnd
rlabel metal1 511 -522 576 -515 5 drain
rlabel metal1 523 -980 588 -973 5 drain
rlabel metal1 518 -1069 588 -1061 1 Gnd
rlabel metal1 351 -1066 421 -1058 1 Gnd
rlabel metal1 356 -977 421 -970 5 drain
rlabel metal1 838 -980 903 -973 5 drain
rlabel metal1 833 -1069 903 -1061 1 Gnd
rlabel metal1 666 -1066 736 -1058 1 Gnd
rlabel metal1 671 -977 736 -970 5 drain
rlabel metal1 224 -1730 289 -1723 5 drain
rlabel metal1 219 -1819 289 -1811 1 Gnd
rlabel metal1 52 -1816 122 -1808 1 Gnd
rlabel metal1 57 -1727 122 -1720 5 drain
rlabel metal1 703 -1384 768 -1377 5 drain
rlabel metal1 698 -1473 768 -1465 1 Gnd
rlabel metal1 865 -1476 935 -1468 1 Gnd
rlabel metal1 870 -1387 935 -1380 5 drain
rlabel metal1 388 -1384 453 -1377 5 drain
rlabel metal1 383 -1473 453 -1465 1 Gnd
rlabel metal1 550 -1476 620 -1468 1 Gnd
rlabel metal1 555 -1387 620 -1380 5 drain
rlabel metal1 273 -1793 281 -1769 1 P1
rlabel metal1 1315 -971 1380 -964 5 drain
rlabel metal1 1310 -1060 1380 -1052 1 Gnd
rlabel metal1 1477 -1063 1547 -1055 1 Gnd
rlabel metal1 1482 -974 1547 -967 5 drain
rlabel metal1 1000 -971 1065 -964 5 drain
rlabel metal1 995 -1060 1065 -1052 1 Gnd
rlabel metal1 1162 -1063 1232 -1055 1 Gnd
rlabel metal1 1167 -974 1232 -967 5 drain
rlabel metal1 919 -1450 927 -1426 1 P2
rlabel metal1 690 -519 755 -512 5 drain
rlabel metal1 1531 -1037 1539 -1013 1 P3
rlabel polysilicon 381 183 386 191 1 f3
rlabel polysilicon 385 -350 389 -344 1 f2
rlabel polysilicon 95 184 97 197 1 f4
rlabel metal1 636 -252 638 -239 1 f5
rlabel metal1 732 -413 734 -400 1 f6
rlabel polysilicon 1046 -353 1048 -340 1 f7
rlabel polysilicon 400 -681 400 -663 1 f8
rlabel metal2 621 -731 623 -713 1 f9
rlabel polysilicon 729 -635 731 -617 1 f10
rlabel metal1 1284 -596 1286 -578 1 f11
rlabel polysilicon 317 -1024 324 -1022 1 f12
rlabel polysilicon 725 -1130 728 -1126 1 f13
rlabel metal1 957 -1130 959 -1106 1 f14
rlabel metal1 1042 -1296 1044 -1272 1 f15
rlabel metal1 1300 -1091 1302 -1067 1 f16
rlabel polysilicon 1357 -1220 1360 -1212 1 f17
rlabel metal1 1575 -1185 1578 -1177 7 f18
rlabel polysilicon 745 -1634 748 -1626 1 f19
rlabel polysilicon 67 -149 70 -134 1 A2B3
rlabel polysilicon 112 -264 115 -249 1 A3B2
rlabel metal1 42 -742 45 -727 1 A3B1
rlabel polysilicon 95 -637 98 -622 1 A2B2
rlabel polysilicon 95 -968 98 -953 1 A3B0
rlabel polysilicon 67 -1026 70 -1011 1 A2B1
rlabel polysilicon 67 -1402 70 -1387 1 A2B0
rlabel polysilicon 95 -1467 98 -1452 1 A1B1
rlabel polysilicon 425 -1505 428 -1490 1 A0B2
rlabel polysilicon 66 -1777 69 -1762 1 A1B0
rlabel polysilicon 95 -1845 98 -1830 1 A0B1
rlabel polysilicon 393 -1092 396 -1078 1 A1B2
<< end >>
